magic
tech sky130A
magscale 1 2
timestamp 1623775656
<< obsli1 >>
rect 1104 1309 198812 199563
<< obsm1 >>
rect 198 76 199810 199980
<< metal2 >>
rect 846 199200 902 200000
rect 2502 199200 2558 200000
rect 4250 199200 4306 200000
rect 5998 199200 6054 200000
rect 7746 199200 7802 200000
rect 9494 199200 9550 200000
rect 11242 199200 11298 200000
rect 12990 199200 13046 200000
rect 14738 199200 14794 200000
rect 16486 199200 16542 200000
rect 18234 199200 18290 200000
rect 19890 199200 19946 200000
rect 21638 199200 21694 200000
rect 23386 199200 23442 200000
rect 25134 199200 25190 200000
rect 26882 199200 26938 200000
rect 28630 199200 28686 200000
rect 30378 199200 30434 200000
rect 32126 199200 32182 200000
rect 33874 199200 33930 200000
rect 35622 199200 35678 200000
rect 37278 199200 37334 200000
rect 39026 199200 39082 200000
rect 40774 199200 40830 200000
rect 42522 199200 42578 200000
rect 44270 199200 44326 200000
rect 46018 199200 46074 200000
rect 47766 199200 47822 200000
rect 49514 199200 49570 200000
rect 51262 199200 51318 200000
rect 53010 199200 53066 200000
rect 54758 199200 54814 200000
rect 56414 199200 56470 200000
rect 58162 199200 58218 200000
rect 59910 199200 59966 200000
rect 61658 199200 61714 200000
rect 63406 199200 63462 200000
rect 65154 199200 65210 200000
rect 66902 199200 66958 200000
rect 68650 199200 68706 200000
rect 70398 199200 70454 200000
rect 72146 199200 72202 200000
rect 73802 199200 73858 200000
rect 75550 199200 75606 200000
rect 77298 199200 77354 200000
rect 79046 199200 79102 200000
rect 80794 199200 80850 200000
rect 82542 199200 82598 200000
rect 84290 199200 84346 200000
rect 86038 199200 86094 200000
rect 87786 199200 87842 200000
rect 89534 199200 89590 200000
rect 91282 199200 91338 200000
rect 92938 199200 92994 200000
rect 94686 199200 94742 200000
rect 96434 199200 96490 200000
rect 98182 199200 98238 200000
rect 99930 199200 99986 200000
rect 101678 199200 101734 200000
rect 103426 199200 103482 200000
rect 105174 199200 105230 200000
rect 106922 199200 106978 200000
rect 108670 199200 108726 200000
rect 110326 199200 110382 200000
rect 112074 199200 112130 200000
rect 113822 199200 113878 200000
rect 115570 199200 115626 200000
rect 117318 199200 117374 200000
rect 119066 199200 119122 200000
rect 120814 199200 120870 200000
rect 122562 199200 122618 200000
rect 124310 199200 124366 200000
rect 126058 199200 126114 200000
rect 127806 199200 127862 200000
rect 129462 199200 129518 200000
rect 131210 199200 131266 200000
rect 132958 199200 133014 200000
rect 134706 199200 134762 200000
rect 136454 199200 136510 200000
rect 138202 199200 138258 200000
rect 139950 199200 140006 200000
rect 141698 199200 141754 200000
rect 143446 199200 143502 200000
rect 145194 199200 145250 200000
rect 146850 199200 146906 200000
rect 148598 199200 148654 200000
rect 150346 199200 150402 200000
rect 152094 199200 152150 200000
rect 153842 199200 153898 200000
rect 155590 199200 155646 200000
rect 157338 199200 157394 200000
rect 159086 199200 159142 200000
rect 160834 199200 160890 200000
rect 162582 199200 162638 200000
rect 164330 199200 164386 200000
rect 165986 199200 166042 200000
rect 167734 199200 167790 200000
rect 169482 199200 169538 200000
rect 171230 199200 171286 200000
rect 172978 199200 173034 200000
rect 174726 199200 174782 200000
rect 176474 199200 176530 200000
rect 178222 199200 178278 200000
rect 179970 199200 180026 200000
rect 181718 199200 181774 200000
rect 183374 199200 183430 200000
rect 185122 199200 185178 200000
rect 186870 199200 186926 200000
rect 188618 199200 188674 200000
rect 190366 199200 190422 200000
rect 192114 199200 192170 200000
rect 193862 199200 193918 200000
rect 195610 199200 195666 200000
rect 197358 199200 197414 200000
rect 199106 199200 199162 200000
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26238 0 26294 800
rect 26606 0 26662 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31942 0 31998 800
rect 32310 0 32366 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34794 0 34850 800
rect 35162 0 35218 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41326 0 41382 800
rect 41694 0 41750 800
rect 42154 0 42210 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43350 0 43406 800
rect 43718 0 43774 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45742 0 45798 800
rect 46202 0 46258 800
rect 46570 0 46626 800
rect 47030 0 47086 800
rect 47398 0 47454 800
rect 47858 0 47914 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49882 0 49938 800
rect 50250 0 50306 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52734 0 52790 800
rect 53102 0 53158 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55126 0 55182 800
rect 55586 0 55642 800
rect 55954 0 56010 800
rect 56414 0 56470 800
rect 56782 0 56838 800
rect 57150 0 57206 800
rect 57610 0 57666 800
rect 57978 0 58034 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 60002 0 60058 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61290 0 61346 800
rect 61658 0 61714 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 64142 0 64198 800
rect 64510 0 64566 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65706 0 65762 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66994 0 67050 800
rect 67362 0 67418 800
rect 67730 0 67786 800
rect 68190 0 68246 800
rect 68558 0 68614 800
rect 69018 0 69074 800
rect 69386 0 69442 800
rect 69846 0 69902 800
rect 70214 0 70270 800
rect 70582 0 70638 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71870 0 71926 800
rect 72238 0 72294 800
rect 72698 0 72754 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74722 0 74778 800
rect 75090 0 75146 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76286 0 76342 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77574 0 77630 800
rect 77942 0 77998 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79138 0 79194 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80426 0 80482 800
rect 80794 0 80850 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84106 0 84162 800
rect 84474 0 84530 800
rect 84842 0 84898 800
rect 85302 0 85358 800
rect 85670 0 85726 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86958 0 87014 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 88154 0 88210 800
rect 88522 0 88578 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89810 0 89866 800
rect 90178 0 90234 800
rect 90546 0 90602 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91834 0 91890 800
rect 92202 0 92258 800
rect 92662 0 92718 800
rect 93030 0 93086 800
rect 93398 0 93454 800
rect 93858 0 93914 800
rect 94226 0 94282 800
rect 94686 0 94742 800
rect 95054 0 95110 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97538 0 97594 800
rect 97906 0 97962 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99562 0 99618 800
rect 99930 0 99986 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101954 0 102010 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 104070 0 104126 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 106094 0 106150 800
rect 106462 0 106518 800
rect 106922 0 106978 800
rect 107290 0 107346 800
rect 107658 0 107714 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108946 0 109002 800
rect 109314 0 109370 800
rect 109774 0 109830 800
rect 110142 0 110198 800
rect 110510 0 110566 800
rect 110970 0 111026 800
rect 111338 0 111394 800
rect 111798 0 111854 800
rect 112166 0 112222 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113822 0 113878 800
rect 114190 0 114246 800
rect 114650 0 114706 800
rect 115018 0 115074 800
rect 115478 0 115534 800
rect 115846 0 115902 800
rect 116214 0 116270 800
rect 116674 0 116730 800
rect 117042 0 117098 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118330 0 118386 800
rect 118698 0 118754 800
rect 119066 0 119122 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121918 0 121974 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123206 0 123262 800
rect 123574 0 123630 800
rect 124034 0 124090 800
rect 124402 0 124458 800
rect 124770 0 124826 800
rect 125230 0 125286 800
rect 125598 0 125654 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126886 0 126942 800
rect 127254 0 127310 800
rect 127622 0 127678 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128910 0 128966 800
rect 129278 0 129334 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130934 0 130990 800
rect 131302 0 131358 800
rect 131762 0 131818 800
rect 132130 0 132186 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134614 0 134670 800
rect 134982 0 135038 800
rect 135350 0 135406 800
rect 135810 0 135866 800
rect 136178 0 136234 800
rect 136638 0 136694 800
rect 137006 0 137062 800
rect 137466 0 137522 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138662 0 138718 800
rect 139030 0 139086 800
rect 139490 0 139546 800
rect 139858 0 139914 800
rect 140318 0 140374 800
rect 140686 0 140742 800
rect 141054 0 141110 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 143170 0 143226 800
rect 143538 0 143594 800
rect 143906 0 143962 800
rect 144366 0 144422 800
rect 144734 0 144790 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 146022 0 146078 800
rect 146390 0 146446 800
rect 146758 0 146814 800
rect 147218 0 147274 800
rect 147586 0 147642 800
rect 148046 0 148102 800
rect 148414 0 148470 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149610 0 149666 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150898 0 150954 800
rect 151266 0 151322 800
rect 151726 0 151782 800
rect 152094 0 152150 800
rect 152462 0 152518 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153750 0 153806 800
rect 154118 0 154174 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155314 0 155370 800
rect 155774 0 155830 800
rect 156142 0 156198 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158626 0 158682 800
rect 158994 0 159050 800
rect 159454 0 159510 800
rect 159822 0 159878 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161478 0 161534 800
rect 161846 0 161902 800
rect 162306 0 162362 800
rect 162674 0 162730 800
rect 163134 0 163190 800
rect 163502 0 163558 800
rect 163870 0 163926 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165158 0 165214 800
rect 165526 0 165582 800
rect 165986 0 166042 800
rect 166354 0 166410 800
rect 166722 0 166778 800
rect 167182 0 167238 800
rect 167550 0 167606 800
rect 168010 0 168066 800
rect 168378 0 168434 800
rect 168838 0 168894 800
rect 169206 0 169262 800
rect 169574 0 169630 800
rect 170034 0 170090 800
rect 170402 0 170458 800
rect 170862 0 170918 800
rect 171230 0 171286 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172886 0 172942 800
rect 173254 0 173310 800
rect 173714 0 173770 800
rect 174082 0 174138 800
rect 174542 0 174598 800
rect 174910 0 174966 800
rect 175278 0 175334 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176566 0 176622 800
rect 176934 0 176990 800
rect 177394 0 177450 800
rect 177762 0 177818 800
rect 178130 0 178186 800
rect 178590 0 178646 800
rect 178958 0 179014 800
rect 179418 0 179474 800
rect 179786 0 179842 800
rect 180246 0 180302 800
rect 180614 0 180670 800
rect 180982 0 181038 800
rect 181442 0 181498 800
rect 181810 0 181866 800
rect 182270 0 182326 800
rect 182638 0 182694 800
rect 183098 0 183154 800
rect 183466 0 183522 800
rect 183834 0 183890 800
rect 184294 0 184350 800
rect 184662 0 184718 800
rect 185122 0 185178 800
rect 185490 0 185546 800
rect 185950 0 186006 800
rect 186318 0 186374 800
rect 186686 0 186742 800
rect 187146 0 187202 800
rect 187514 0 187570 800
rect 187974 0 188030 800
rect 188342 0 188398 800
rect 188802 0 188858 800
rect 189170 0 189226 800
rect 189538 0 189594 800
rect 189998 0 190054 800
rect 190366 0 190422 800
rect 190826 0 190882 800
rect 191194 0 191250 800
rect 191654 0 191710 800
rect 192022 0 192078 800
rect 192390 0 192446 800
rect 192850 0 192906 800
rect 193218 0 193274 800
rect 193678 0 193734 800
rect 194046 0 194102 800
rect 194506 0 194562 800
rect 194874 0 194930 800
rect 195242 0 195298 800
rect 195702 0 195758 800
rect 196070 0 196126 800
rect 196530 0 196586 800
rect 196898 0 196954 800
rect 197358 0 197414 800
rect 197726 0 197782 800
rect 198094 0 198150 800
rect 198554 0 198610 800
rect 198922 0 198978 800
rect 199382 0 199438 800
rect 199750 0 199806 800
<< obsm2 >>
rect 204 199144 790 199986
rect 958 199144 2446 199986
rect 2614 199144 4194 199986
rect 4362 199144 5942 199986
rect 6110 199144 7690 199986
rect 7858 199144 9438 199986
rect 9606 199144 11186 199986
rect 11354 199144 12934 199986
rect 13102 199144 14682 199986
rect 14850 199144 16430 199986
rect 16598 199144 18178 199986
rect 18346 199144 19834 199986
rect 20002 199144 21582 199986
rect 21750 199144 23330 199986
rect 23498 199144 25078 199986
rect 25246 199144 26826 199986
rect 26994 199144 28574 199986
rect 28742 199144 30322 199986
rect 30490 199144 32070 199986
rect 32238 199144 33818 199986
rect 33986 199144 35566 199986
rect 35734 199144 37222 199986
rect 37390 199144 38970 199986
rect 39138 199144 40718 199986
rect 40886 199144 42466 199986
rect 42634 199144 44214 199986
rect 44382 199144 45962 199986
rect 46130 199144 47710 199986
rect 47878 199144 49458 199986
rect 49626 199144 51206 199986
rect 51374 199144 52954 199986
rect 53122 199144 54702 199986
rect 54870 199144 56358 199986
rect 56526 199144 58106 199986
rect 58274 199144 59854 199986
rect 60022 199144 61602 199986
rect 61770 199144 63350 199986
rect 63518 199144 65098 199986
rect 65266 199144 66846 199986
rect 67014 199144 68594 199986
rect 68762 199144 70342 199986
rect 70510 199144 72090 199986
rect 72258 199144 73746 199986
rect 73914 199144 75494 199986
rect 75662 199144 77242 199986
rect 77410 199144 78990 199986
rect 79158 199144 80738 199986
rect 80906 199144 82486 199986
rect 82654 199144 84234 199986
rect 84402 199144 85982 199986
rect 86150 199144 87730 199986
rect 87898 199144 89478 199986
rect 89646 199144 91226 199986
rect 91394 199144 92882 199986
rect 93050 199144 94630 199986
rect 94798 199144 96378 199986
rect 96546 199144 98126 199986
rect 98294 199144 99874 199986
rect 100042 199144 101622 199986
rect 101790 199144 103370 199986
rect 103538 199144 105118 199986
rect 105286 199144 106866 199986
rect 107034 199144 108614 199986
rect 108782 199144 110270 199986
rect 110438 199144 112018 199986
rect 112186 199144 113766 199986
rect 113934 199144 115514 199986
rect 115682 199144 117262 199986
rect 117430 199144 119010 199986
rect 119178 199144 120758 199986
rect 120926 199144 122506 199986
rect 122674 199144 124254 199986
rect 124422 199144 126002 199986
rect 126170 199144 127750 199986
rect 127918 199144 129406 199986
rect 129574 199144 131154 199986
rect 131322 199144 132902 199986
rect 133070 199144 134650 199986
rect 134818 199144 136398 199986
rect 136566 199144 138146 199986
rect 138314 199144 139894 199986
rect 140062 199144 141642 199986
rect 141810 199144 143390 199986
rect 143558 199144 145138 199986
rect 145306 199144 146794 199986
rect 146962 199144 148542 199986
rect 148710 199144 150290 199986
rect 150458 199144 152038 199986
rect 152206 199144 153786 199986
rect 153954 199144 155534 199986
rect 155702 199144 157282 199986
rect 157450 199144 159030 199986
rect 159198 199144 160778 199986
rect 160946 199144 162526 199986
rect 162694 199144 164274 199986
rect 164442 199144 165930 199986
rect 166098 199144 167678 199986
rect 167846 199144 169426 199986
rect 169594 199144 171174 199986
rect 171342 199144 172922 199986
rect 173090 199144 174670 199986
rect 174838 199144 176418 199986
rect 176586 199144 178166 199986
rect 178334 199144 179914 199986
rect 180082 199144 181662 199986
rect 181830 199144 183318 199986
rect 183486 199144 185066 199986
rect 185234 199144 186814 199986
rect 186982 199144 188562 199986
rect 188730 199144 190310 199986
rect 190478 199144 192058 199986
rect 192226 199144 193806 199986
rect 193974 199144 195554 199986
rect 195722 199144 197302 199986
rect 197470 199144 199050 199986
rect 199218 199144 199804 199986
rect 204 856 199804 199144
rect 314 70 514 856
rect 682 70 882 856
rect 1050 70 1342 856
rect 1510 70 1710 856
rect 1878 70 2170 856
rect 2338 70 2538 856
rect 2706 70 2906 856
rect 3074 70 3366 856
rect 3534 70 3734 856
rect 3902 70 4194 856
rect 4362 70 4562 856
rect 4730 70 5022 856
rect 5190 70 5390 856
rect 5558 70 5758 856
rect 5926 70 6218 856
rect 6386 70 6586 856
rect 6754 70 7046 856
rect 7214 70 7414 856
rect 7582 70 7874 856
rect 8042 70 8242 856
rect 8410 70 8610 856
rect 8778 70 9070 856
rect 9238 70 9438 856
rect 9606 70 9898 856
rect 10066 70 10266 856
rect 10434 70 10726 856
rect 10894 70 11094 856
rect 11262 70 11462 856
rect 11630 70 11922 856
rect 12090 70 12290 856
rect 12458 70 12750 856
rect 12918 70 13118 856
rect 13286 70 13578 856
rect 13746 70 13946 856
rect 14114 70 14314 856
rect 14482 70 14774 856
rect 14942 70 15142 856
rect 15310 70 15602 856
rect 15770 70 15970 856
rect 16138 70 16430 856
rect 16598 70 16798 856
rect 16966 70 17166 856
rect 17334 70 17626 856
rect 17794 70 17994 856
rect 18162 70 18454 856
rect 18622 70 18822 856
rect 18990 70 19282 856
rect 19450 70 19650 856
rect 19818 70 20018 856
rect 20186 70 20478 856
rect 20646 70 20846 856
rect 21014 70 21306 856
rect 21474 70 21674 856
rect 21842 70 22134 856
rect 22302 70 22502 856
rect 22670 70 22870 856
rect 23038 70 23330 856
rect 23498 70 23698 856
rect 23866 70 24158 856
rect 24326 70 24526 856
rect 24694 70 24986 856
rect 25154 70 25354 856
rect 25522 70 25722 856
rect 25890 70 26182 856
rect 26350 70 26550 856
rect 26718 70 27010 856
rect 27178 70 27378 856
rect 27546 70 27838 856
rect 28006 70 28206 856
rect 28374 70 28574 856
rect 28742 70 29034 856
rect 29202 70 29402 856
rect 29570 70 29862 856
rect 30030 70 30230 856
rect 30398 70 30690 856
rect 30858 70 31058 856
rect 31226 70 31426 856
rect 31594 70 31886 856
rect 32054 70 32254 856
rect 32422 70 32714 856
rect 32882 70 33082 856
rect 33250 70 33542 856
rect 33710 70 33910 856
rect 34078 70 34278 856
rect 34446 70 34738 856
rect 34906 70 35106 856
rect 35274 70 35566 856
rect 35734 70 35934 856
rect 36102 70 36394 856
rect 36562 70 36762 856
rect 36930 70 37130 856
rect 37298 70 37590 856
rect 37758 70 37958 856
rect 38126 70 38418 856
rect 38586 70 38786 856
rect 38954 70 39246 856
rect 39414 70 39614 856
rect 39782 70 39982 856
rect 40150 70 40442 856
rect 40610 70 40810 856
rect 40978 70 41270 856
rect 41438 70 41638 856
rect 41806 70 42098 856
rect 42266 70 42466 856
rect 42634 70 42834 856
rect 43002 70 43294 856
rect 43462 70 43662 856
rect 43830 70 44122 856
rect 44290 70 44490 856
rect 44658 70 44950 856
rect 45118 70 45318 856
rect 45486 70 45686 856
rect 45854 70 46146 856
rect 46314 70 46514 856
rect 46682 70 46974 856
rect 47142 70 47342 856
rect 47510 70 47802 856
rect 47970 70 48170 856
rect 48338 70 48538 856
rect 48706 70 48998 856
rect 49166 70 49366 856
rect 49534 70 49826 856
rect 49994 70 50194 856
rect 50362 70 50654 856
rect 50822 70 51022 856
rect 51190 70 51390 856
rect 51558 70 51850 856
rect 52018 70 52218 856
rect 52386 70 52678 856
rect 52846 70 53046 856
rect 53214 70 53506 856
rect 53674 70 53874 856
rect 54042 70 54242 856
rect 54410 70 54702 856
rect 54870 70 55070 856
rect 55238 70 55530 856
rect 55698 70 55898 856
rect 56066 70 56358 856
rect 56526 70 56726 856
rect 56894 70 57094 856
rect 57262 70 57554 856
rect 57722 70 57922 856
rect 58090 70 58382 856
rect 58550 70 58750 856
rect 58918 70 59210 856
rect 59378 70 59578 856
rect 59746 70 59946 856
rect 60114 70 60406 856
rect 60574 70 60774 856
rect 60942 70 61234 856
rect 61402 70 61602 856
rect 61770 70 62062 856
rect 62230 70 62430 856
rect 62598 70 62798 856
rect 62966 70 63258 856
rect 63426 70 63626 856
rect 63794 70 64086 856
rect 64254 70 64454 856
rect 64622 70 64914 856
rect 65082 70 65282 856
rect 65450 70 65650 856
rect 65818 70 66110 856
rect 66278 70 66478 856
rect 66646 70 66938 856
rect 67106 70 67306 856
rect 67474 70 67674 856
rect 67842 70 68134 856
rect 68302 70 68502 856
rect 68670 70 68962 856
rect 69130 70 69330 856
rect 69498 70 69790 856
rect 69958 70 70158 856
rect 70326 70 70526 856
rect 70694 70 70986 856
rect 71154 70 71354 856
rect 71522 70 71814 856
rect 71982 70 72182 856
rect 72350 70 72642 856
rect 72810 70 73010 856
rect 73178 70 73378 856
rect 73546 70 73838 856
rect 74006 70 74206 856
rect 74374 70 74666 856
rect 74834 70 75034 856
rect 75202 70 75494 856
rect 75662 70 75862 856
rect 76030 70 76230 856
rect 76398 70 76690 856
rect 76858 70 77058 856
rect 77226 70 77518 856
rect 77686 70 77886 856
rect 78054 70 78346 856
rect 78514 70 78714 856
rect 78882 70 79082 856
rect 79250 70 79542 856
rect 79710 70 79910 856
rect 80078 70 80370 856
rect 80538 70 80738 856
rect 80906 70 81198 856
rect 81366 70 81566 856
rect 81734 70 81934 856
rect 82102 70 82394 856
rect 82562 70 82762 856
rect 82930 70 83222 856
rect 83390 70 83590 856
rect 83758 70 84050 856
rect 84218 70 84418 856
rect 84586 70 84786 856
rect 84954 70 85246 856
rect 85414 70 85614 856
rect 85782 70 86074 856
rect 86242 70 86442 856
rect 86610 70 86902 856
rect 87070 70 87270 856
rect 87438 70 87638 856
rect 87806 70 88098 856
rect 88266 70 88466 856
rect 88634 70 88926 856
rect 89094 70 89294 856
rect 89462 70 89754 856
rect 89922 70 90122 856
rect 90290 70 90490 856
rect 90658 70 90950 856
rect 91118 70 91318 856
rect 91486 70 91778 856
rect 91946 70 92146 856
rect 92314 70 92606 856
rect 92774 70 92974 856
rect 93142 70 93342 856
rect 93510 70 93802 856
rect 93970 70 94170 856
rect 94338 70 94630 856
rect 94798 70 94998 856
rect 95166 70 95458 856
rect 95626 70 95826 856
rect 95994 70 96194 856
rect 96362 70 96654 856
rect 96822 70 97022 856
rect 97190 70 97482 856
rect 97650 70 97850 856
rect 98018 70 98310 856
rect 98478 70 98678 856
rect 98846 70 99046 856
rect 99214 70 99506 856
rect 99674 70 99874 856
rect 100042 70 100334 856
rect 100502 70 100702 856
rect 100870 70 101162 856
rect 101330 70 101530 856
rect 101698 70 101898 856
rect 102066 70 102358 856
rect 102526 70 102726 856
rect 102894 70 103186 856
rect 103354 70 103554 856
rect 103722 70 104014 856
rect 104182 70 104382 856
rect 104550 70 104750 856
rect 104918 70 105210 856
rect 105378 70 105578 856
rect 105746 70 106038 856
rect 106206 70 106406 856
rect 106574 70 106866 856
rect 107034 70 107234 856
rect 107402 70 107602 856
rect 107770 70 108062 856
rect 108230 70 108430 856
rect 108598 70 108890 856
rect 109058 70 109258 856
rect 109426 70 109718 856
rect 109886 70 110086 856
rect 110254 70 110454 856
rect 110622 70 110914 856
rect 111082 70 111282 856
rect 111450 70 111742 856
rect 111910 70 112110 856
rect 112278 70 112570 856
rect 112738 70 112938 856
rect 113106 70 113306 856
rect 113474 70 113766 856
rect 113934 70 114134 856
rect 114302 70 114594 856
rect 114762 70 114962 856
rect 115130 70 115422 856
rect 115590 70 115790 856
rect 115958 70 116158 856
rect 116326 70 116618 856
rect 116786 70 116986 856
rect 117154 70 117446 856
rect 117614 70 117814 856
rect 117982 70 118274 856
rect 118442 70 118642 856
rect 118810 70 119010 856
rect 119178 70 119470 856
rect 119638 70 119838 856
rect 120006 70 120298 856
rect 120466 70 120666 856
rect 120834 70 121126 856
rect 121294 70 121494 856
rect 121662 70 121862 856
rect 122030 70 122322 856
rect 122490 70 122690 856
rect 122858 70 123150 856
rect 123318 70 123518 856
rect 123686 70 123978 856
rect 124146 70 124346 856
rect 124514 70 124714 856
rect 124882 70 125174 856
rect 125342 70 125542 856
rect 125710 70 126002 856
rect 126170 70 126370 856
rect 126538 70 126830 856
rect 126998 70 127198 856
rect 127366 70 127566 856
rect 127734 70 128026 856
rect 128194 70 128394 856
rect 128562 70 128854 856
rect 129022 70 129222 856
rect 129390 70 129682 856
rect 129850 70 130050 856
rect 130218 70 130418 856
rect 130586 70 130878 856
rect 131046 70 131246 856
rect 131414 70 131706 856
rect 131874 70 132074 856
rect 132242 70 132534 856
rect 132702 70 132902 856
rect 133070 70 133270 856
rect 133438 70 133730 856
rect 133898 70 134098 856
rect 134266 70 134558 856
rect 134726 70 134926 856
rect 135094 70 135294 856
rect 135462 70 135754 856
rect 135922 70 136122 856
rect 136290 70 136582 856
rect 136750 70 136950 856
rect 137118 70 137410 856
rect 137578 70 137778 856
rect 137946 70 138146 856
rect 138314 70 138606 856
rect 138774 70 138974 856
rect 139142 70 139434 856
rect 139602 70 139802 856
rect 139970 70 140262 856
rect 140430 70 140630 856
rect 140798 70 140998 856
rect 141166 70 141458 856
rect 141626 70 141826 856
rect 141994 70 142286 856
rect 142454 70 142654 856
rect 142822 70 143114 856
rect 143282 70 143482 856
rect 143650 70 143850 856
rect 144018 70 144310 856
rect 144478 70 144678 856
rect 144846 70 145138 856
rect 145306 70 145506 856
rect 145674 70 145966 856
rect 146134 70 146334 856
rect 146502 70 146702 856
rect 146870 70 147162 856
rect 147330 70 147530 856
rect 147698 70 147990 856
rect 148158 70 148358 856
rect 148526 70 148818 856
rect 148986 70 149186 856
rect 149354 70 149554 856
rect 149722 70 150014 856
rect 150182 70 150382 856
rect 150550 70 150842 856
rect 151010 70 151210 856
rect 151378 70 151670 856
rect 151838 70 152038 856
rect 152206 70 152406 856
rect 152574 70 152866 856
rect 153034 70 153234 856
rect 153402 70 153694 856
rect 153862 70 154062 856
rect 154230 70 154522 856
rect 154690 70 154890 856
rect 155058 70 155258 856
rect 155426 70 155718 856
rect 155886 70 156086 856
rect 156254 70 156546 856
rect 156714 70 156914 856
rect 157082 70 157374 856
rect 157542 70 157742 856
rect 157910 70 158110 856
rect 158278 70 158570 856
rect 158738 70 158938 856
rect 159106 70 159398 856
rect 159566 70 159766 856
rect 159934 70 160226 856
rect 160394 70 160594 856
rect 160762 70 160962 856
rect 161130 70 161422 856
rect 161590 70 161790 856
rect 161958 70 162250 856
rect 162418 70 162618 856
rect 162786 70 163078 856
rect 163246 70 163446 856
rect 163614 70 163814 856
rect 163982 70 164274 856
rect 164442 70 164642 856
rect 164810 70 165102 856
rect 165270 70 165470 856
rect 165638 70 165930 856
rect 166098 70 166298 856
rect 166466 70 166666 856
rect 166834 70 167126 856
rect 167294 70 167494 856
rect 167662 70 167954 856
rect 168122 70 168322 856
rect 168490 70 168782 856
rect 168950 70 169150 856
rect 169318 70 169518 856
rect 169686 70 169978 856
rect 170146 70 170346 856
rect 170514 70 170806 856
rect 170974 70 171174 856
rect 171342 70 171634 856
rect 171802 70 172002 856
rect 172170 70 172370 856
rect 172538 70 172830 856
rect 172998 70 173198 856
rect 173366 70 173658 856
rect 173826 70 174026 856
rect 174194 70 174486 856
rect 174654 70 174854 856
rect 175022 70 175222 856
rect 175390 70 175682 856
rect 175850 70 176050 856
rect 176218 70 176510 856
rect 176678 70 176878 856
rect 177046 70 177338 856
rect 177506 70 177706 856
rect 177874 70 178074 856
rect 178242 70 178534 856
rect 178702 70 178902 856
rect 179070 70 179362 856
rect 179530 70 179730 856
rect 179898 70 180190 856
rect 180358 70 180558 856
rect 180726 70 180926 856
rect 181094 70 181386 856
rect 181554 70 181754 856
rect 181922 70 182214 856
rect 182382 70 182582 856
rect 182750 70 183042 856
rect 183210 70 183410 856
rect 183578 70 183778 856
rect 183946 70 184238 856
rect 184406 70 184606 856
rect 184774 70 185066 856
rect 185234 70 185434 856
rect 185602 70 185894 856
rect 186062 70 186262 856
rect 186430 70 186630 856
rect 186798 70 187090 856
rect 187258 70 187458 856
rect 187626 70 187918 856
rect 188086 70 188286 856
rect 188454 70 188746 856
rect 188914 70 189114 856
rect 189282 70 189482 856
rect 189650 70 189942 856
rect 190110 70 190310 856
rect 190478 70 190770 856
rect 190938 70 191138 856
rect 191306 70 191598 856
rect 191766 70 191966 856
rect 192134 70 192334 856
rect 192502 70 192794 856
rect 192962 70 193162 856
rect 193330 70 193622 856
rect 193790 70 193990 856
rect 194158 70 194450 856
rect 194618 70 194818 856
rect 194986 70 195186 856
rect 195354 70 195646 856
rect 195814 70 196014 856
rect 196182 70 196474 856
rect 196642 70 196842 856
rect 197010 70 197302 856
rect 197470 70 197670 856
rect 197838 70 198038 856
rect 198206 70 198498 856
rect 198666 70 198866 856
rect 199034 70 199326 856
rect 199494 70 199694 856
<< metal3 >>
rect 0 99968 800 100088
<< obsm3 >>
rect 800 100168 188848 198661
rect 880 99888 188848 100168
rect 800 171 188848 99888
<< metal4 >>
rect 4208 2128 4528 197520
rect 4868 2176 5188 197472
rect 5528 2176 5848 197472
rect 6188 2176 6508 197472
rect 19568 2128 19888 197520
rect 20228 2176 20548 197472
rect 20888 2176 21208 197472
rect 21548 2176 21868 197472
rect 34928 2128 35248 197520
rect 35588 2176 35908 197472
rect 36248 2176 36568 197472
rect 36908 2176 37228 197472
rect 50288 2128 50608 197520
rect 50948 2176 51268 197472
rect 51608 2176 51928 197472
rect 52268 2176 52588 197472
rect 65648 2128 65968 197520
rect 66308 2176 66628 197472
rect 66968 2176 67288 197472
rect 67628 2176 67948 197472
rect 81008 2128 81328 197520
rect 81668 2176 81988 197472
rect 82328 2176 82648 197472
rect 82988 2176 83308 197472
rect 96368 2128 96688 197520
rect 97028 2176 97348 197472
rect 97688 2176 98008 197472
rect 98348 2176 98668 197472
rect 111728 2128 112048 197520
rect 112388 2176 112708 197472
rect 113048 2176 113368 197472
rect 113708 2176 114028 197472
rect 127088 2128 127408 197520
rect 127748 2176 128068 197472
rect 128408 2176 128728 197472
rect 129068 2176 129388 197472
rect 142448 2128 142768 197520
rect 143108 2176 143428 197472
rect 143768 2176 144088 197472
rect 144428 2176 144748 197472
rect 157808 2128 158128 197520
rect 158468 2176 158788 197472
rect 159128 2176 159448 197472
rect 159788 2176 160108 197472
rect 173168 2128 173488 197520
rect 173828 2176 174148 197472
rect 174488 2176 174808 197472
rect 175148 2176 175468 197472
rect 188528 2128 188848 197520
rect 189188 2176 189508 197472
rect 189848 2176 190168 197472
rect 190508 2176 190828 197472
<< obsm4 >>
rect 3187 197600 184309 198661
rect 3187 2048 4128 197600
rect 4608 197552 19488 197600
rect 4608 2096 4788 197552
rect 5268 2096 5448 197552
rect 5928 2096 6108 197552
rect 6588 2096 19488 197552
rect 19968 197552 34848 197600
rect 4608 2048 19488 2096
rect 19968 2096 20148 197552
rect 20628 2096 20808 197552
rect 21288 2096 21468 197552
rect 21948 2096 34848 197552
rect 35328 197552 50208 197600
rect 19968 2048 34848 2096
rect 35328 2096 35508 197552
rect 35988 2096 36168 197552
rect 36648 2096 36828 197552
rect 37308 2096 50208 197552
rect 50688 197552 65568 197600
rect 35328 2048 50208 2096
rect 50688 2096 50868 197552
rect 51348 2096 51528 197552
rect 52008 2096 52188 197552
rect 52668 2096 65568 197552
rect 66048 197552 80928 197600
rect 50688 2048 65568 2096
rect 66048 2096 66228 197552
rect 66708 2096 66888 197552
rect 67368 2096 67548 197552
rect 68028 2096 80928 197552
rect 81408 197552 96288 197600
rect 66048 2048 80928 2096
rect 81408 2096 81588 197552
rect 82068 2096 82248 197552
rect 82728 2096 82908 197552
rect 83388 2096 96288 197552
rect 96768 197552 111648 197600
rect 81408 2048 96288 2096
rect 96768 2096 96948 197552
rect 97428 2096 97608 197552
rect 98088 2096 98268 197552
rect 98748 2096 111648 197552
rect 112128 197552 127008 197600
rect 96768 2048 111648 2096
rect 112128 2096 112308 197552
rect 112788 2096 112968 197552
rect 113448 2096 113628 197552
rect 114108 2096 127008 197552
rect 127488 197552 142368 197600
rect 112128 2048 127008 2096
rect 127488 2096 127668 197552
rect 128148 2096 128328 197552
rect 128808 2096 128988 197552
rect 129468 2096 142368 197552
rect 142848 197552 157728 197600
rect 127488 2048 142368 2096
rect 142848 2096 143028 197552
rect 143508 2096 143688 197552
rect 144168 2096 144348 197552
rect 144828 2096 157728 197552
rect 158208 197552 173088 197600
rect 142848 2048 157728 2096
rect 158208 2096 158388 197552
rect 158868 2096 159048 197552
rect 159528 2096 159708 197552
rect 160188 2096 173088 197552
rect 173568 197552 184309 197600
rect 158208 2048 173088 2096
rect 173568 2096 173748 197552
rect 174228 2096 174408 197552
rect 174888 2096 175068 197552
rect 175548 2096 184309 197552
rect 173568 2048 184309 2096
rect 3187 902 184309 2048
<< obsm5 >>
rect 30476 860 153892 197020
<< labels >>
rlabel metal2 s 846 199200 902 200000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 53010 199200 53066 200000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 58162 199200 58218 200000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 63406 199200 63462 200000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 68650 199200 68706 200000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 73802 199200 73858 200000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 79046 199200 79102 200000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 84290 199200 84346 200000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 89534 199200 89590 200000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 94686 199200 94742 200000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 99930 199200 99986 200000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5998 199200 6054 200000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 105174 199200 105230 200000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 110326 199200 110382 200000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 115570 199200 115626 200000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 120814 199200 120870 200000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 126058 199200 126114 200000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 131210 199200 131266 200000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 136454 199200 136510 200000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 141698 199200 141754 200000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 146850 199200 146906 200000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 152094 199200 152150 200000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 11242 199200 11298 200000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 157338 199200 157394 200000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 162582 199200 162638 200000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 167734 199200 167790 200000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 172978 199200 173034 200000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 178222 199200 178278 200000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 183374 199200 183430 200000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 188618 199200 188674 200000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 193862 199200 193918 200000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 16486 199200 16542 200000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 21638 199200 21694 200000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 26882 199200 26938 200000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 32126 199200 32182 200000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 37278 199200 37334 200000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 42522 199200 42578 200000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 47766 199200 47822 200000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2502 199200 2558 200000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 54758 199200 54814 200000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 59910 199200 59966 200000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 65154 199200 65210 200000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 70398 199200 70454 200000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 75550 199200 75606 200000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 80794 199200 80850 200000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 86038 199200 86094 200000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 91282 199200 91338 200000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 96434 199200 96490 200000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 101678 199200 101734 200000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7746 199200 7802 200000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 106922 199200 106978 200000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 112074 199200 112130 200000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 117318 199200 117374 200000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 122562 199200 122618 200000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 127806 199200 127862 200000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 132958 199200 133014 200000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 138202 199200 138258 200000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 143446 199200 143502 200000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 148598 199200 148654 200000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 153842 199200 153898 200000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 12990 199200 13046 200000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 159086 199200 159142 200000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 164330 199200 164386 200000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 169482 199200 169538 200000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 174726 199200 174782 200000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 179970 199200 180026 200000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 185122 199200 185178 200000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 190366 199200 190422 200000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 195610 199200 195666 200000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 18234 199200 18290 200000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 23386 199200 23442 200000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 28630 199200 28686 200000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 33874 199200 33930 200000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 39026 199200 39082 200000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 44270 199200 44326 200000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 49514 199200 49570 200000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4250 199200 4306 200000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 56414 199200 56470 200000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 61658 199200 61714 200000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 66902 199200 66958 200000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 72146 199200 72202 200000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 77298 199200 77354 200000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 82542 199200 82598 200000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 87786 199200 87842 200000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 92938 199200 92994 200000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 98182 199200 98238 200000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 103426 199200 103482 200000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 9494 199200 9550 200000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 108670 199200 108726 200000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 113822 199200 113878 200000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 119066 199200 119122 200000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 124310 199200 124366 200000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 129462 199200 129518 200000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 134706 199200 134762 200000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 139950 199200 140006 200000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 145194 199200 145250 200000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 150346 199200 150402 200000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 155590 199200 155646 200000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 14738 199200 14794 200000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 160834 199200 160890 200000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 165986 199200 166042 200000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 171230 199200 171286 200000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 176474 199200 176530 200000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 181718 199200 181774 200000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 186870 199200 186926 200000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 192114 199200 192170 200000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 197358 199200 197414 200000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 19890 199200 19946 200000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 25134 199200 25190 200000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 30378 199200 30434 200000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 35622 199200 35678 200000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 40774 199200 40830 200000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 46018 199200 46074 200000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 51262 199200 51318 200000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 199750 0 199806 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 199106 199200 199162 200000 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 176566 0 176622 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 180246 0 180302 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 181442 0 181498 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 185122 0 185178 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 187514 0 187570 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 192390 0 192446 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 194874 0 194930 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 155774 0 155830 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 165986 0 166042 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 167182 0 167238 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 169574 0 169630 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 174542 0 174598 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 176934 0 176990 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 178130 0 178186 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 179418 0 179474 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 180614 0 180670 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 181810 0 181866 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 183098 0 183154 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 184294 0 184350 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 186686 0 186742 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 187974 0 188030 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 189170 0 189226 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 190366 0 190422 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 191654 0 191710 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 192850 0 192906 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 194046 0 194102 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 195242 0 195298 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 196530 0 196586 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 197726 0 197782 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 198922 0 198978 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 131762 0 131818 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 135350 0 135406 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 139030 0 139086 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 142710 0 142766 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 143906 0 143962 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 145194 0 145250 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 146390 0 146446 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 151266 0 151322 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 154946 0 155002 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 158626 0 158682 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 159822 0 159878 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 161018 0 161074 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 163502 0 163558 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 164698 0 164754 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 174910 0 174966 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 177394 0 177450 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 179786 0 179842 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 184662 0 184718 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 193218 0 193274 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 195702 0 195758 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 199382 0 199438 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 615 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 189188 2176 189508 197472 6 vccd2
port 621 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 197472 6 vccd2
port 622 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 197472 6 vccd2
port 623 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 197472 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 197472 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 197472 6 vccd2
port 626 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 197472 6 vccd2
port 627 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 197472 6 vssd2
port 628 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 197472 6 vssd2
port 629 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 197472 6 vssd2
port 630 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 197472 6 vssd2
port 631 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 197472 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 197472 6 vssd2
port 633 nsew ground bidirectional
rlabel metal4 s 189848 2176 190168 197472 6 vdda1
port 634 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 197472 6 vdda1
port 635 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 197472 6 vdda1
port 636 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 197472 6 vdda1
port 637 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 197472 6 vdda1
port 638 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 197472 6 vdda1
port 639 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 197472 6 vdda1
port 640 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 197472 6 vssa1
port 641 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 197472 6 vssa1
port 642 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 197472 6 vssa1
port 643 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 197472 6 vssa1
port 644 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 197472 6 vssa1
port 645 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 197472 6 vssa1
port 646 nsew ground bidirectional
rlabel metal4 s 190508 2176 190828 197472 6 vdda2
port 647 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 197472 6 vdda2
port 648 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 197472 6 vdda2
port 649 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 197472 6 vdda2
port 650 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 197472 6 vdda2
port 651 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 197472 6 vdda2
port 652 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 197472 6 vdda2
port 653 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 197472 6 vssa2
port 654 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 197472 6 vssa2
port 655 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 197472 6 vssa2
port 656 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 197472 6 vssa2
port 657 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 197472 6 vssa2
port 658 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 197472 6 vssa2
port 659 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 200000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 112474510
string GDS_START 1258184
<< end >>

