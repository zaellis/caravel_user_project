// File name:   CAN_receiver.sv
// Created:     12/1/2020
// Author:      Zachary Ellis
// Version:     2.0  Integration into full controller
// Description: Top module of CAN receiver project

module CAN_receiver (
    input clk,
    input nRST,
    input [3:0] TS1,
    input [3:0] TS2,
    input CANRX,
    input tx_busy,
    input [1:0] error_state,
    input fifo_clear,
    input enable_overrun,
    input [19:0] mask_enable,
    input [30:0] filter_0, //this is a yosys thing since you cant do input [31:0] [19:0]
    input [30:0] mask_0,
    input [30:0] filter_1,
    input [30:0] mask_1,
    input [30:0] filter_2,
    input [30:0] mask_2,
    input [30:0] filter_3,
    input [30:0] mask_3,
    input [30:0] filter_4,
    input [30:0] mask_4,
    input [30:0] filter_5,
    input [30:0] mask_5,
    input [30:0] filter_6,
    input [30:0] mask_6,
    input [30:0] filter_7,
    input [30:0] mask_7,
    input [30:0] filter_8,
    input [30:0] mask_8,
    input [30:0] filter_9,
    input [30:0] mask_9,
    input [30:0] filter_10,
    input [30:0] mask_10,
    input [30:0] filter_11,
    input [30:0] mask_11,
    input [30:0] filter_12,
    input [30:0] mask_12,
    input [30:0] filter_13,
    input [30:0] mask_13,
    input [30:0] filter_14,
    input [30:0] mask_14,
    input [30:0] filter_15,
    input [30:0] mask_15,
    input [30:0] filter_16,
    input [30:0] mask_16,
    input [30:0] filter_17,
    input [30:0] mask_17,
    input [30:0] filter_18,
    input [30:0] mask_18,
    input [30:0] filter_19,
    input [30:0] mask_19,
    input read_fifo,
    output ACK,
    output busy,
    output bitstuff_error,
    output form_error,
    output [1:0] rx_err_code,
    output CRC_Error,
    output bitstrobe,
    output tx_strobe,
    output curr_sample,
    output [3:0] occupancy,
    output full,
    output empty,
    output overrun,
    output [31:0] data_L,
    output [31:0] data_H,
    output [28:0] ID_out,
    output [3:0] pkt_size_out,
    output RTR_out,
    output EXT_out,
    output [4:0] fmi_out,
    output fifo_read
);

    wire SOF, bitstuff, dataphase, end_data, load_byte, endCRC, edgedet;
    wire [3:0] pkt_size, byte_num, byte_select;
    wire [7:0] payload;
    wire [28:0] CAN_ID;
    wire stopCRC;
    wire RTR, EXT;
    wire pkt_done, new_ID;

    edgedetect U1 (
        .clk(clk),
        .nRST(nRST),
        .CANRX(CANRX),
        .edgedet(edgedet)
    );

    timer U2 (
        .clk(clk),
        .nRST(nRST),
        .TS1(TS1),
        .TS2(TS2),
        .edgedet(edgedet),
        .bitstuff(bitstuff),
        .dataphase(dataphase),
        .pkt_size(pkt_size),
        .bitstrobe(bitstrobe),
        .tx_strobe(tx_strobe),
        .byte_complete(load_byte),
        .byte_num(byte_num),
        .end_data(end_data)
    );

    CRCcheck U3 (
        .clk(clk),
        .bitstrobe(bitstrobe),
        .tx_strobe(tx_strobe),
        .endCRC(endCRC),
        .stopCRC(stopCRC),
        .nRST(nRST),
        .bitstuff(bitstuff),
        .pkt_size(pkt_size),
        .SOF(SOF),
        .CANRX(CANRX),
        .ACK(ACK),
        .CRCerror(CRC_Error)
    );

    RCU U4 (
        .clk(clk),
        .bitstrobe(bitstrobe),
        .nRST(nRST),
        .CANRX(CANRX),
        .tx_busy(tx_busy),
        .error_state(error_state),
        .CRC_err(CRC_Error),
        .enddata(end_data),
        .endCRC(endCRC),
        .stopCRC(stopCRC),
        .busy(busy),
        .Dataphase(dataphase),
        .bitstuff(bitstuff),
        .bitstuff_error(bitstuff_error),
        .form_error(form_error),
        .rx_err_code(rx_err_code),
        .pkt_size(pkt_size),
        .msg_id(CAN_ID),
        .payload(payload),
        .RTR(RTR),
        .EXT(EXT),
        .curr_sample(curr_sample),
        .SOF(SOF),
        .pkt_done(pkt_done),
        .new_ID(new_ID)
    );

    fifo U5 (
        .clk(clk),
        .nRST(nRST),
        .clear(fifo_clear),
        .ID(CAN_ID),
        .data(payload),
        .data_index(byte_num),
        .load_data(load_byte),
        .pkt_size(pkt_size),
        .RTR(RTR),
        .EXT(EXT),
        .pkt_done(pkt_done),
        .enable_overrun(enable_overrun),
        .new_ID(new_ID),
        .mask_enable(mask_enable),
        .filter_0(filter_0),
        .mask_0(mask_0),
        .filter_1(filter_1),
        .mask_1(mask_1),
        .filter_2(filter_2),
        .mask_2(mask_2),
        .filter_3(filter_3),
        .mask_3(mask_3),
        .filter_4(filter_4),
        .mask_4(mask_4),
        .filter_5(filter_5),
        .mask_5(mask_5),
        .filter_6(filter_6),
        .mask_6(mask_6),
        .filter_7(filter_7),
        .mask_7(mask_7),
        .filter_8(filter_8),
        .mask_8(mask_8),
        .filter_9(filter_9),
        .mask_9(mask_9),
        .filter_10(filter_10),
        .mask_10(mask_10),
        .filter_11(filter_11),
        .mask_11(mask_11),
        .filter_12(filter_12),
        .mask_12(mask_12),
        .filter_13(filter_13),
        .mask_13(mask_13),
        .filter_14(filter_14),
        .mask_14(mask_14),
        .filter_15(filter_15),
        .mask_15(mask_15),
        .filter_16(filter_16),
        .mask_16(mask_16),
        .filter_17(filter_17),
        .mask_17(mask_17),
        .filter_18(filter_18),
        .mask_18(mask_18),
        .filter_19(filter_19),
        .mask_19(mask_19),
        .read_fifo(read_fifo),
        .occupancy(occupancy),
        .full(full),
        .empty(empty),
        .overrun(overrun),
        .data_L(data_L),
        .data_H(data_H),
        .ID_out(ID_out),
        .pkt_size_out(pkt_size_out),
        .RTR_out(RTR_out),
        .EXT_out(EXT_out),
        .fmi_out(fmi_out),
        .fifo_read(fifo_read)
    );    

endmodule