magic
tech sky130A
magscale 1 2
timestamp 1624577832
<< obsli1 >>
rect 29 2159 338836 337841
<< obsm1 >>
rect 14 1912 339650 337872
<< metal2 >>
rect 1490 339200 1546 340000
rect 4434 339200 4490 340000
rect 7378 339200 7434 340000
rect 10322 339200 10378 340000
rect 13266 339200 13322 340000
rect 16210 339200 16266 340000
rect 19154 339200 19210 340000
rect 22098 339200 22154 340000
rect 25134 339200 25190 340000
rect 28078 339200 28134 340000
rect 31022 339200 31078 340000
rect 33966 339200 34022 340000
rect 36910 339200 36966 340000
rect 39854 339200 39910 340000
rect 42798 339200 42854 340000
rect 45834 339200 45890 340000
rect 48778 339200 48834 340000
rect 51722 339200 51778 340000
rect 54666 339200 54722 340000
rect 57610 339200 57666 340000
rect 60554 339200 60610 340000
rect 63498 339200 63554 340000
rect 66534 339200 66590 340000
rect 69478 339200 69534 340000
rect 72422 339200 72478 340000
rect 75366 339200 75422 340000
rect 78310 339200 78366 340000
rect 81254 339200 81310 340000
rect 84198 339200 84254 340000
rect 87234 339200 87290 340000
rect 90178 339200 90234 340000
rect 93122 339200 93178 340000
rect 96066 339200 96122 340000
rect 99010 339200 99066 340000
rect 101954 339200 102010 340000
rect 104898 339200 104954 340000
rect 107934 339200 107990 340000
rect 110878 339200 110934 340000
rect 113822 339200 113878 340000
rect 116766 339200 116822 340000
rect 119710 339200 119766 340000
rect 122654 339200 122710 340000
rect 125598 339200 125654 340000
rect 128542 339200 128598 340000
rect 131578 339200 131634 340000
rect 134522 339200 134578 340000
rect 137466 339200 137522 340000
rect 140410 339200 140466 340000
rect 143354 339200 143410 340000
rect 146298 339200 146354 340000
rect 149242 339200 149298 340000
rect 152278 339200 152334 340000
rect 155222 339200 155278 340000
rect 158166 339200 158222 340000
rect 161110 339200 161166 340000
rect 164054 339200 164110 340000
rect 166998 339200 167054 340000
rect 169942 339200 169998 340000
rect 172978 339200 173034 340000
rect 175922 339200 175978 340000
rect 178866 339200 178922 340000
rect 181810 339200 181866 340000
rect 184754 339200 184810 340000
rect 187698 339200 187754 340000
rect 190642 339200 190698 340000
rect 193678 339200 193734 340000
rect 196622 339200 196678 340000
rect 199566 339200 199622 340000
rect 202510 339200 202566 340000
rect 205454 339200 205510 340000
rect 208398 339200 208454 340000
rect 211342 339200 211398 340000
rect 214378 339200 214434 340000
rect 217322 339200 217378 340000
rect 220266 339200 220322 340000
rect 223210 339200 223266 340000
rect 226154 339200 226210 340000
rect 229098 339200 229154 340000
rect 232042 339200 232098 340000
rect 234986 339200 235042 340000
rect 238022 339200 238078 340000
rect 240966 339200 241022 340000
rect 243910 339200 243966 340000
rect 246854 339200 246910 340000
rect 249798 339200 249854 340000
rect 252742 339200 252798 340000
rect 255686 339200 255742 340000
rect 258722 339200 258778 340000
rect 261666 339200 261722 340000
rect 264610 339200 264666 340000
rect 267554 339200 267610 340000
rect 270498 339200 270554 340000
rect 273442 339200 273498 340000
rect 276386 339200 276442 340000
rect 279422 339200 279478 340000
rect 282366 339200 282422 340000
rect 285310 339200 285366 340000
rect 288254 339200 288310 340000
rect 291198 339200 291254 340000
rect 294142 339200 294198 340000
rect 297086 339200 297142 340000
rect 300122 339200 300178 340000
rect 303066 339200 303122 340000
rect 306010 339200 306066 340000
rect 308954 339200 309010 340000
rect 311898 339200 311954 340000
rect 314842 339200 314898 340000
rect 317786 339200 317842 340000
rect 320822 339200 320878 340000
rect 323766 339200 323822 340000
rect 326710 339200 326766 340000
rect 329654 339200 329710 340000
rect 332598 339200 332654 340000
rect 335542 339200 335598 340000
rect 338486 339200 338542 340000
rect 294 0 350 800
rect 938 0 994 800
rect 1674 0 1730 800
rect 2318 0 2374 800
rect 3054 0 3110 800
rect 3698 0 3754 800
rect 4434 0 4490 800
rect 5078 0 5134 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7838 0 7894 800
rect 8574 0 8630 800
rect 9218 0 9274 800
rect 9954 0 10010 800
rect 10598 0 10654 800
rect 11334 0 11390 800
rect 11978 0 12034 800
rect 12714 0 12770 800
rect 13450 0 13506 800
rect 14094 0 14150 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16210 0 16266 800
rect 16854 0 16910 800
rect 17590 0 17646 800
rect 18234 0 18290 800
rect 18970 0 19026 800
rect 19614 0 19670 800
rect 20350 0 20406 800
rect 20994 0 21050 800
rect 21730 0 21786 800
rect 22374 0 22430 800
rect 23110 0 23166 800
rect 23754 0 23810 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25870 0 25926 800
rect 26606 0 26662 800
rect 27250 0 27306 800
rect 27986 0 28042 800
rect 28630 0 28686 800
rect 29366 0 29422 800
rect 30010 0 30066 800
rect 30746 0 30802 800
rect 31390 0 31446 800
rect 32126 0 32182 800
rect 32770 0 32826 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34886 0 34942 800
rect 35530 0 35586 800
rect 36266 0 36322 800
rect 36910 0 36966 800
rect 37646 0 37702 800
rect 38382 0 38438 800
rect 39026 0 39082 800
rect 39762 0 39818 800
rect 40406 0 40462 800
rect 41142 0 41198 800
rect 41786 0 41842 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43902 0 43958 800
rect 44546 0 44602 800
rect 45282 0 45338 800
rect 45926 0 45982 800
rect 46662 0 46718 800
rect 47306 0 47362 800
rect 48042 0 48098 800
rect 48686 0 48742 800
rect 49422 0 49478 800
rect 50066 0 50122 800
rect 50802 0 50858 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 52918 0 52974 800
rect 53562 0 53618 800
rect 54298 0 54354 800
rect 54942 0 54998 800
rect 55678 0 55734 800
rect 56322 0 56378 800
rect 57058 0 57114 800
rect 57702 0 57758 800
rect 58438 0 58494 800
rect 59082 0 59138 800
rect 59818 0 59874 800
rect 60462 0 60518 800
rect 61198 0 61254 800
rect 61842 0 61898 800
rect 62578 0 62634 800
rect 63314 0 63370 800
rect 63958 0 64014 800
rect 64694 0 64750 800
rect 65338 0 65394 800
rect 66074 0 66130 800
rect 66718 0 66774 800
rect 67454 0 67510 800
rect 68098 0 68154 800
rect 68834 0 68890 800
rect 69478 0 69534 800
rect 70214 0 70270 800
rect 70858 0 70914 800
rect 71594 0 71650 800
rect 72238 0 72294 800
rect 72974 0 73030 800
rect 73618 0 73674 800
rect 74354 0 74410 800
rect 74998 0 75054 800
rect 75734 0 75790 800
rect 76470 0 76526 800
rect 77114 0 77170 800
rect 77850 0 77906 800
rect 78494 0 78550 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 80610 0 80666 800
rect 81254 0 81310 800
rect 81990 0 82046 800
rect 82634 0 82690 800
rect 83370 0 83426 800
rect 84014 0 84070 800
rect 84750 0 84806 800
rect 85394 0 85450 800
rect 86130 0 86186 800
rect 86774 0 86830 800
rect 87510 0 87566 800
rect 88154 0 88210 800
rect 88890 0 88946 800
rect 89626 0 89682 800
rect 90270 0 90326 800
rect 91006 0 91062 800
rect 91650 0 91706 800
rect 92386 0 92442 800
rect 93030 0 93086 800
rect 93766 0 93822 800
rect 94410 0 94466 800
rect 95146 0 95202 800
rect 95790 0 95846 800
rect 96526 0 96582 800
rect 97170 0 97226 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99286 0 99342 800
rect 99930 0 99986 800
rect 100666 0 100722 800
rect 101402 0 101458 800
rect 102046 0 102102 800
rect 102782 0 102838 800
rect 103426 0 103482 800
rect 104162 0 104218 800
rect 104806 0 104862 800
rect 105542 0 105598 800
rect 106186 0 106242 800
rect 106922 0 106978 800
rect 107566 0 107622 800
rect 108302 0 108358 800
rect 108946 0 109002 800
rect 109682 0 109738 800
rect 110326 0 110382 800
rect 111062 0 111118 800
rect 111706 0 111762 800
rect 112442 0 112498 800
rect 113086 0 113142 800
rect 113822 0 113878 800
rect 114558 0 114614 800
rect 115202 0 115258 800
rect 115938 0 115994 800
rect 116582 0 116638 800
rect 117318 0 117374 800
rect 117962 0 118018 800
rect 118698 0 118754 800
rect 119342 0 119398 800
rect 120078 0 120134 800
rect 120722 0 120778 800
rect 121458 0 121514 800
rect 122102 0 122158 800
rect 122838 0 122894 800
rect 123482 0 123538 800
rect 124218 0 124274 800
rect 124862 0 124918 800
rect 125598 0 125654 800
rect 126334 0 126390 800
rect 126978 0 127034 800
rect 127714 0 127770 800
rect 128358 0 128414 800
rect 129094 0 129150 800
rect 129738 0 129794 800
rect 130474 0 130530 800
rect 131118 0 131174 800
rect 131854 0 131910 800
rect 132498 0 132554 800
rect 133234 0 133290 800
rect 133878 0 133934 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 135994 0 136050 800
rect 136638 0 136694 800
rect 137374 0 137430 800
rect 138018 0 138074 800
rect 138754 0 138810 800
rect 139490 0 139546 800
rect 140134 0 140190 800
rect 140870 0 140926 800
rect 141514 0 141570 800
rect 142250 0 142306 800
rect 142894 0 142950 800
rect 143630 0 143686 800
rect 144274 0 144330 800
rect 145010 0 145066 800
rect 145654 0 145710 800
rect 146390 0 146446 800
rect 147034 0 147090 800
rect 147770 0 147826 800
rect 148414 0 148470 800
rect 149150 0 149206 800
rect 149794 0 149850 800
rect 150530 0 150586 800
rect 151174 0 151230 800
rect 151910 0 151966 800
rect 152646 0 152702 800
rect 153290 0 153346 800
rect 154026 0 154082 800
rect 154670 0 154726 800
rect 155406 0 155462 800
rect 156050 0 156106 800
rect 156786 0 156842 800
rect 157430 0 157486 800
rect 158166 0 158222 800
rect 158810 0 158866 800
rect 159546 0 159602 800
rect 160190 0 160246 800
rect 160926 0 160982 800
rect 161570 0 161626 800
rect 162306 0 162362 800
rect 162950 0 163006 800
rect 163686 0 163742 800
rect 164422 0 164478 800
rect 165066 0 165122 800
rect 165802 0 165858 800
rect 166446 0 166502 800
rect 167182 0 167238 800
rect 167826 0 167882 800
rect 168562 0 168618 800
rect 169206 0 169262 800
rect 169942 0 169998 800
rect 170586 0 170642 800
rect 171322 0 171378 800
rect 171966 0 172022 800
rect 172702 0 172758 800
rect 173346 0 173402 800
rect 174082 0 174138 800
rect 174726 0 174782 800
rect 175462 0 175518 800
rect 176106 0 176162 800
rect 176842 0 176898 800
rect 177578 0 177634 800
rect 178222 0 178278 800
rect 178958 0 179014 800
rect 179602 0 179658 800
rect 180338 0 180394 800
rect 180982 0 181038 800
rect 181718 0 181774 800
rect 182362 0 182418 800
rect 183098 0 183154 800
rect 183742 0 183798 800
rect 184478 0 184534 800
rect 185122 0 185178 800
rect 185858 0 185914 800
rect 186502 0 186558 800
rect 187238 0 187294 800
rect 187882 0 187938 800
rect 188618 0 188674 800
rect 189354 0 189410 800
rect 189998 0 190054 800
rect 190734 0 190790 800
rect 191378 0 191434 800
rect 192114 0 192170 800
rect 192758 0 192814 800
rect 193494 0 193550 800
rect 194138 0 194194 800
rect 194874 0 194930 800
rect 195518 0 195574 800
rect 196254 0 196310 800
rect 196898 0 196954 800
rect 197634 0 197690 800
rect 198278 0 198334 800
rect 199014 0 199070 800
rect 199658 0 199714 800
rect 200394 0 200450 800
rect 201038 0 201094 800
rect 201774 0 201830 800
rect 202510 0 202566 800
rect 203154 0 203210 800
rect 203890 0 203946 800
rect 204534 0 204590 800
rect 205270 0 205326 800
rect 205914 0 205970 800
rect 206650 0 206706 800
rect 207294 0 207350 800
rect 208030 0 208086 800
rect 208674 0 208730 800
rect 209410 0 209466 800
rect 210054 0 210110 800
rect 210790 0 210846 800
rect 211434 0 211490 800
rect 212170 0 212226 800
rect 212814 0 212870 800
rect 213550 0 213606 800
rect 214194 0 214250 800
rect 214930 0 214986 800
rect 215666 0 215722 800
rect 216310 0 216366 800
rect 217046 0 217102 800
rect 217690 0 217746 800
rect 218426 0 218482 800
rect 219070 0 219126 800
rect 219806 0 219862 800
rect 220450 0 220506 800
rect 221186 0 221242 800
rect 221830 0 221886 800
rect 222566 0 222622 800
rect 223210 0 223266 800
rect 223946 0 224002 800
rect 224590 0 224646 800
rect 225326 0 225382 800
rect 225970 0 226026 800
rect 226706 0 226762 800
rect 227442 0 227498 800
rect 228086 0 228142 800
rect 228822 0 228878 800
rect 229466 0 229522 800
rect 230202 0 230258 800
rect 230846 0 230902 800
rect 231582 0 231638 800
rect 232226 0 232282 800
rect 232962 0 233018 800
rect 233606 0 233662 800
rect 234342 0 234398 800
rect 234986 0 235042 800
rect 235722 0 235778 800
rect 236366 0 236422 800
rect 237102 0 237158 800
rect 237746 0 237802 800
rect 238482 0 238538 800
rect 239126 0 239182 800
rect 239862 0 239918 800
rect 240598 0 240654 800
rect 241242 0 241298 800
rect 241978 0 242034 800
rect 242622 0 242678 800
rect 243358 0 243414 800
rect 244002 0 244058 800
rect 244738 0 244794 800
rect 245382 0 245438 800
rect 246118 0 246174 800
rect 246762 0 246818 800
rect 247498 0 247554 800
rect 248142 0 248198 800
rect 248878 0 248934 800
rect 249522 0 249578 800
rect 250258 0 250314 800
rect 250902 0 250958 800
rect 251638 0 251694 800
rect 252374 0 252430 800
rect 253018 0 253074 800
rect 253754 0 253810 800
rect 254398 0 254454 800
rect 255134 0 255190 800
rect 255778 0 255834 800
rect 256514 0 256570 800
rect 257158 0 257214 800
rect 257894 0 257950 800
rect 258538 0 258594 800
rect 259274 0 259330 800
rect 259918 0 259974 800
rect 260654 0 260710 800
rect 261298 0 261354 800
rect 262034 0 262090 800
rect 262678 0 262734 800
rect 263414 0 263470 800
rect 264058 0 264114 800
rect 264794 0 264850 800
rect 265530 0 265586 800
rect 266174 0 266230 800
rect 266910 0 266966 800
rect 267554 0 267610 800
rect 268290 0 268346 800
rect 268934 0 268990 800
rect 269670 0 269726 800
rect 270314 0 270370 800
rect 271050 0 271106 800
rect 271694 0 271750 800
rect 272430 0 272486 800
rect 273074 0 273130 800
rect 273810 0 273866 800
rect 274454 0 274510 800
rect 275190 0 275246 800
rect 275834 0 275890 800
rect 276570 0 276626 800
rect 277214 0 277270 800
rect 277950 0 278006 800
rect 278686 0 278742 800
rect 279330 0 279386 800
rect 280066 0 280122 800
rect 280710 0 280766 800
rect 281446 0 281502 800
rect 282090 0 282146 800
rect 282826 0 282882 800
rect 283470 0 283526 800
rect 284206 0 284262 800
rect 284850 0 284906 800
rect 285586 0 285642 800
rect 286230 0 286286 800
rect 286966 0 287022 800
rect 287610 0 287666 800
rect 288346 0 288402 800
rect 288990 0 289046 800
rect 289726 0 289782 800
rect 290462 0 290518 800
rect 291106 0 291162 800
rect 291842 0 291898 800
rect 292486 0 292542 800
rect 293222 0 293278 800
rect 293866 0 293922 800
rect 294602 0 294658 800
rect 295246 0 295302 800
rect 295982 0 296038 800
rect 296626 0 296682 800
rect 297362 0 297418 800
rect 298006 0 298062 800
rect 298742 0 298798 800
rect 299386 0 299442 800
rect 300122 0 300178 800
rect 300766 0 300822 800
rect 301502 0 301558 800
rect 302146 0 302202 800
rect 302882 0 302938 800
rect 303618 0 303674 800
rect 304262 0 304318 800
rect 304998 0 305054 800
rect 305642 0 305698 800
rect 306378 0 306434 800
rect 307022 0 307078 800
rect 307758 0 307814 800
rect 308402 0 308458 800
rect 309138 0 309194 800
rect 309782 0 309838 800
rect 310518 0 310574 800
rect 311162 0 311218 800
rect 311898 0 311954 800
rect 312542 0 312598 800
rect 313278 0 313334 800
rect 313922 0 313978 800
rect 314658 0 314714 800
rect 315394 0 315450 800
rect 316038 0 316094 800
rect 316774 0 316830 800
rect 317418 0 317474 800
rect 318154 0 318210 800
rect 318798 0 318854 800
rect 319534 0 319590 800
rect 320178 0 320234 800
rect 320914 0 320970 800
rect 321558 0 321614 800
rect 322294 0 322350 800
rect 322938 0 322994 800
rect 323674 0 323730 800
rect 324318 0 324374 800
rect 325054 0 325110 800
rect 325698 0 325754 800
rect 326434 0 326490 800
rect 327078 0 327134 800
rect 327814 0 327870 800
rect 328550 0 328606 800
rect 329194 0 329250 800
rect 329930 0 329986 800
rect 330574 0 330630 800
rect 331310 0 331366 800
rect 331954 0 332010 800
rect 332690 0 332746 800
rect 333334 0 333390 800
rect 334070 0 334126 800
rect 334714 0 334770 800
rect 335450 0 335506 800
rect 336094 0 336150 800
rect 336830 0 336886 800
rect 337474 0 337530 800
rect 338210 0 338266 800
rect 338854 0 338910 800
rect 339590 0 339646 800
<< obsm2 >>
rect 18 339144 1434 339200
rect 1602 339144 4378 339200
rect 4546 339144 7322 339200
rect 7490 339144 10266 339200
rect 10434 339144 13210 339200
rect 13378 339144 16154 339200
rect 16322 339144 19098 339200
rect 19266 339144 22042 339200
rect 22210 339144 25078 339200
rect 25246 339144 28022 339200
rect 28190 339144 30966 339200
rect 31134 339144 33910 339200
rect 34078 339144 36854 339200
rect 37022 339144 39798 339200
rect 39966 339144 42742 339200
rect 42910 339144 45778 339200
rect 45946 339144 48722 339200
rect 48890 339144 51666 339200
rect 51834 339144 54610 339200
rect 54778 339144 57554 339200
rect 57722 339144 60498 339200
rect 60666 339144 63442 339200
rect 63610 339144 66478 339200
rect 66646 339144 69422 339200
rect 69590 339144 72366 339200
rect 72534 339144 75310 339200
rect 75478 339144 78254 339200
rect 78422 339144 81198 339200
rect 81366 339144 84142 339200
rect 84310 339144 87178 339200
rect 87346 339144 90122 339200
rect 90290 339144 93066 339200
rect 93234 339144 96010 339200
rect 96178 339144 98954 339200
rect 99122 339144 101898 339200
rect 102066 339144 104842 339200
rect 105010 339144 107878 339200
rect 108046 339144 110822 339200
rect 110990 339144 113766 339200
rect 113934 339144 116710 339200
rect 116878 339144 119654 339200
rect 119822 339144 122598 339200
rect 122766 339144 125542 339200
rect 125710 339144 128486 339200
rect 128654 339144 131522 339200
rect 131690 339144 134466 339200
rect 134634 339144 137410 339200
rect 137578 339144 140354 339200
rect 140522 339144 143298 339200
rect 143466 339144 146242 339200
rect 146410 339144 149186 339200
rect 149354 339144 152222 339200
rect 152390 339144 155166 339200
rect 155334 339144 158110 339200
rect 158278 339144 161054 339200
rect 161222 339144 163998 339200
rect 164166 339144 166942 339200
rect 167110 339144 169886 339200
rect 170054 339144 172922 339200
rect 173090 339144 175866 339200
rect 176034 339144 178810 339200
rect 178978 339144 181754 339200
rect 181922 339144 184698 339200
rect 184866 339144 187642 339200
rect 187810 339144 190586 339200
rect 190754 339144 193622 339200
rect 193790 339144 196566 339200
rect 196734 339144 199510 339200
rect 199678 339144 202454 339200
rect 202622 339144 205398 339200
rect 205566 339144 208342 339200
rect 208510 339144 211286 339200
rect 211454 339144 214322 339200
rect 214490 339144 217266 339200
rect 217434 339144 220210 339200
rect 220378 339144 223154 339200
rect 223322 339144 226098 339200
rect 226266 339144 229042 339200
rect 229210 339144 231986 339200
rect 232154 339144 234930 339200
rect 235098 339144 237966 339200
rect 238134 339144 240910 339200
rect 241078 339144 243854 339200
rect 244022 339144 246798 339200
rect 246966 339144 249742 339200
rect 249910 339144 252686 339200
rect 252854 339144 255630 339200
rect 255798 339144 258666 339200
rect 258834 339144 261610 339200
rect 261778 339144 264554 339200
rect 264722 339144 267498 339200
rect 267666 339144 270442 339200
rect 270610 339144 273386 339200
rect 273554 339144 276330 339200
rect 276498 339144 279366 339200
rect 279534 339144 282310 339200
rect 282478 339144 285254 339200
rect 285422 339144 288198 339200
rect 288366 339144 291142 339200
rect 291310 339144 294086 339200
rect 294254 339144 297030 339200
rect 297198 339144 300066 339200
rect 300234 339144 303010 339200
rect 303178 339144 305954 339200
rect 306122 339144 308898 339200
rect 309066 339144 311842 339200
rect 312010 339144 314786 339200
rect 314954 339144 317730 339200
rect 317898 339144 320766 339200
rect 320934 339144 323710 339200
rect 323878 339144 326654 339200
rect 326822 339144 329598 339200
rect 329766 339144 332542 339200
rect 332710 339144 335486 339200
rect 335654 339144 338430 339200
rect 338598 339144 339644 339200
rect 18 856 339644 339144
rect 18 800 238 856
rect 406 800 882 856
rect 1050 800 1618 856
rect 1786 800 2262 856
rect 2430 800 2998 856
rect 3166 800 3642 856
rect 3810 800 4378 856
rect 4546 800 5022 856
rect 5190 800 5758 856
rect 5926 800 6402 856
rect 6570 800 7138 856
rect 7306 800 7782 856
rect 7950 800 8518 856
rect 8686 800 9162 856
rect 9330 800 9898 856
rect 10066 800 10542 856
rect 10710 800 11278 856
rect 11446 800 11922 856
rect 12090 800 12658 856
rect 12826 800 13394 856
rect 13562 800 14038 856
rect 14206 800 14774 856
rect 14942 800 15418 856
rect 15586 800 16154 856
rect 16322 800 16798 856
rect 16966 800 17534 856
rect 17702 800 18178 856
rect 18346 800 18914 856
rect 19082 800 19558 856
rect 19726 800 20294 856
rect 20462 800 20938 856
rect 21106 800 21674 856
rect 21842 800 22318 856
rect 22486 800 23054 856
rect 23222 800 23698 856
rect 23866 800 24434 856
rect 24602 800 25078 856
rect 25246 800 25814 856
rect 25982 800 26550 856
rect 26718 800 27194 856
rect 27362 800 27930 856
rect 28098 800 28574 856
rect 28742 800 29310 856
rect 29478 800 29954 856
rect 30122 800 30690 856
rect 30858 800 31334 856
rect 31502 800 32070 856
rect 32238 800 32714 856
rect 32882 800 33450 856
rect 33618 800 34094 856
rect 34262 800 34830 856
rect 34998 800 35474 856
rect 35642 800 36210 856
rect 36378 800 36854 856
rect 37022 800 37590 856
rect 37758 800 38326 856
rect 38494 800 38970 856
rect 39138 800 39706 856
rect 39874 800 40350 856
rect 40518 800 41086 856
rect 41254 800 41730 856
rect 41898 800 42466 856
rect 42634 800 43110 856
rect 43278 800 43846 856
rect 44014 800 44490 856
rect 44658 800 45226 856
rect 45394 800 45870 856
rect 46038 800 46606 856
rect 46774 800 47250 856
rect 47418 800 47986 856
rect 48154 800 48630 856
rect 48798 800 49366 856
rect 49534 800 50010 856
rect 50178 800 50746 856
rect 50914 800 51482 856
rect 51650 800 52126 856
rect 52294 800 52862 856
rect 53030 800 53506 856
rect 53674 800 54242 856
rect 54410 800 54886 856
rect 55054 800 55622 856
rect 55790 800 56266 856
rect 56434 800 57002 856
rect 57170 800 57646 856
rect 57814 800 58382 856
rect 58550 800 59026 856
rect 59194 800 59762 856
rect 59930 800 60406 856
rect 60574 800 61142 856
rect 61310 800 61786 856
rect 61954 800 62522 856
rect 62690 800 63258 856
rect 63426 800 63902 856
rect 64070 800 64638 856
rect 64806 800 65282 856
rect 65450 800 66018 856
rect 66186 800 66662 856
rect 66830 800 67398 856
rect 67566 800 68042 856
rect 68210 800 68778 856
rect 68946 800 69422 856
rect 69590 800 70158 856
rect 70326 800 70802 856
rect 70970 800 71538 856
rect 71706 800 72182 856
rect 72350 800 72918 856
rect 73086 800 73562 856
rect 73730 800 74298 856
rect 74466 800 74942 856
rect 75110 800 75678 856
rect 75846 800 76414 856
rect 76582 800 77058 856
rect 77226 800 77794 856
rect 77962 800 78438 856
rect 78606 800 79174 856
rect 79342 800 79818 856
rect 79986 800 80554 856
rect 80722 800 81198 856
rect 81366 800 81934 856
rect 82102 800 82578 856
rect 82746 800 83314 856
rect 83482 800 83958 856
rect 84126 800 84694 856
rect 84862 800 85338 856
rect 85506 800 86074 856
rect 86242 800 86718 856
rect 86886 800 87454 856
rect 87622 800 88098 856
rect 88266 800 88834 856
rect 89002 800 89570 856
rect 89738 800 90214 856
rect 90382 800 90950 856
rect 91118 800 91594 856
rect 91762 800 92330 856
rect 92498 800 92974 856
rect 93142 800 93710 856
rect 93878 800 94354 856
rect 94522 800 95090 856
rect 95258 800 95734 856
rect 95902 800 96470 856
rect 96638 800 97114 856
rect 97282 800 97850 856
rect 98018 800 98494 856
rect 98662 800 99230 856
rect 99398 800 99874 856
rect 100042 800 100610 856
rect 100778 800 101346 856
rect 101514 800 101990 856
rect 102158 800 102726 856
rect 102894 800 103370 856
rect 103538 800 104106 856
rect 104274 800 104750 856
rect 104918 800 105486 856
rect 105654 800 106130 856
rect 106298 800 106866 856
rect 107034 800 107510 856
rect 107678 800 108246 856
rect 108414 800 108890 856
rect 109058 800 109626 856
rect 109794 800 110270 856
rect 110438 800 111006 856
rect 111174 800 111650 856
rect 111818 800 112386 856
rect 112554 800 113030 856
rect 113198 800 113766 856
rect 113934 800 114502 856
rect 114670 800 115146 856
rect 115314 800 115882 856
rect 116050 800 116526 856
rect 116694 800 117262 856
rect 117430 800 117906 856
rect 118074 800 118642 856
rect 118810 800 119286 856
rect 119454 800 120022 856
rect 120190 800 120666 856
rect 120834 800 121402 856
rect 121570 800 122046 856
rect 122214 800 122782 856
rect 122950 800 123426 856
rect 123594 800 124162 856
rect 124330 800 124806 856
rect 124974 800 125542 856
rect 125710 800 126278 856
rect 126446 800 126922 856
rect 127090 800 127658 856
rect 127826 800 128302 856
rect 128470 800 129038 856
rect 129206 800 129682 856
rect 129850 800 130418 856
rect 130586 800 131062 856
rect 131230 800 131798 856
rect 131966 800 132442 856
rect 132610 800 133178 856
rect 133346 800 133822 856
rect 133990 800 134558 856
rect 134726 800 135202 856
rect 135370 800 135938 856
rect 136106 800 136582 856
rect 136750 800 137318 856
rect 137486 800 137962 856
rect 138130 800 138698 856
rect 138866 800 139434 856
rect 139602 800 140078 856
rect 140246 800 140814 856
rect 140982 800 141458 856
rect 141626 800 142194 856
rect 142362 800 142838 856
rect 143006 800 143574 856
rect 143742 800 144218 856
rect 144386 800 144954 856
rect 145122 800 145598 856
rect 145766 800 146334 856
rect 146502 800 146978 856
rect 147146 800 147714 856
rect 147882 800 148358 856
rect 148526 800 149094 856
rect 149262 800 149738 856
rect 149906 800 150474 856
rect 150642 800 151118 856
rect 151286 800 151854 856
rect 152022 800 152590 856
rect 152758 800 153234 856
rect 153402 800 153970 856
rect 154138 800 154614 856
rect 154782 800 155350 856
rect 155518 800 155994 856
rect 156162 800 156730 856
rect 156898 800 157374 856
rect 157542 800 158110 856
rect 158278 800 158754 856
rect 158922 800 159490 856
rect 159658 800 160134 856
rect 160302 800 160870 856
rect 161038 800 161514 856
rect 161682 800 162250 856
rect 162418 800 162894 856
rect 163062 800 163630 856
rect 163798 800 164366 856
rect 164534 800 165010 856
rect 165178 800 165746 856
rect 165914 800 166390 856
rect 166558 800 167126 856
rect 167294 800 167770 856
rect 167938 800 168506 856
rect 168674 800 169150 856
rect 169318 800 169886 856
rect 170054 800 170530 856
rect 170698 800 171266 856
rect 171434 800 171910 856
rect 172078 800 172646 856
rect 172814 800 173290 856
rect 173458 800 174026 856
rect 174194 800 174670 856
rect 174838 800 175406 856
rect 175574 800 176050 856
rect 176218 800 176786 856
rect 176954 800 177522 856
rect 177690 800 178166 856
rect 178334 800 178902 856
rect 179070 800 179546 856
rect 179714 800 180282 856
rect 180450 800 180926 856
rect 181094 800 181662 856
rect 181830 800 182306 856
rect 182474 800 183042 856
rect 183210 800 183686 856
rect 183854 800 184422 856
rect 184590 800 185066 856
rect 185234 800 185802 856
rect 185970 800 186446 856
rect 186614 800 187182 856
rect 187350 800 187826 856
rect 187994 800 188562 856
rect 188730 800 189298 856
rect 189466 800 189942 856
rect 190110 800 190678 856
rect 190846 800 191322 856
rect 191490 800 192058 856
rect 192226 800 192702 856
rect 192870 800 193438 856
rect 193606 800 194082 856
rect 194250 800 194818 856
rect 194986 800 195462 856
rect 195630 800 196198 856
rect 196366 800 196842 856
rect 197010 800 197578 856
rect 197746 800 198222 856
rect 198390 800 198958 856
rect 199126 800 199602 856
rect 199770 800 200338 856
rect 200506 800 200982 856
rect 201150 800 201718 856
rect 201886 800 202454 856
rect 202622 800 203098 856
rect 203266 800 203834 856
rect 204002 800 204478 856
rect 204646 800 205214 856
rect 205382 800 205858 856
rect 206026 800 206594 856
rect 206762 800 207238 856
rect 207406 800 207974 856
rect 208142 800 208618 856
rect 208786 800 209354 856
rect 209522 800 209998 856
rect 210166 800 210734 856
rect 210902 800 211378 856
rect 211546 800 212114 856
rect 212282 800 212758 856
rect 212926 800 213494 856
rect 213662 800 214138 856
rect 214306 800 214874 856
rect 215042 800 215610 856
rect 215778 800 216254 856
rect 216422 800 216990 856
rect 217158 800 217634 856
rect 217802 800 218370 856
rect 218538 800 219014 856
rect 219182 800 219750 856
rect 219918 800 220394 856
rect 220562 800 221130 856
rect 221298 800 221774 856
rect 221942 800 222510 856
rect 222678 800 223154 856
rect 223322 800 223890 856
rect 224058 800 224534 856
rect 224702 800 225270 856
rect 225438 800 225914 856
rect 226082 800 226650 856
rect 226818 800 227386 856
rect 227554 800 228030 856
rect 228198 800 228766 856
rect 228934 800 229410 856
rect 229578 800 230146 856
rect 230314 800 230790 856
rect 230958 800 231526 856
rect 231694 800 232170 856
rect 232338 800 232906 856
rect 233074 800 233550 856
rect 233718 800 234286 856
rect 234454 800 234930 856
rect 235098 800 235666 856
rect 235834 800 236310 856
rect 236478 800 237046 856
rect 237214 800 237690 856
rect 237858 800 238426 856
rect 238594 800 239070 856
rect 239238 800 239806 856
rect 239974 800 240542 856
rect 240710 800 241186 856
rect 241354 800 241922 856
rect 242090 800 242566 856
rect 242734 800 243302 856
rect 243470 800 243946 856
rect 244114 800 244682 856
rect 244850 800 245326 856
rect 245494 800 246062 856
rect 246230 800 246706 856
rect 246874 800 247442 856
rect 247610 800 248086 856
rect 248254 800 248822 856
rect 248990 800 249466 856
rect 249634 800 250202 856
rect 250370 800 250846 856
rect 251014 800 251582 856
rect 251750 800 252318 856
rect 252486 800 252962 856
rect 253130 800 253698 856
rect 253866 800 254342 856
rect 254510 800 255078 856
rect 255246 800 255722 856
rect 255890 800 256458 856
rect 256626 800 257102 856
rect 257270 800 257838 856
rect 258006 800 258482 856
rect 258650 800 259218 856
rect 259386 800 259862 856
rect 260030 800 260598 856
rect 260766 800 261242 856
rect 261410 800 261978 856
rect 262146 800 262622 856
rect 262790 800 263358 856
rect 263526 800 264002 856
rect 264170 800 264738 856
rect 264906 800 265474 856
rect 265642 800 266118 856
rect 266286 800 266854 856
rect 267022 800 267498 856
rect 267666 800 268234 856
rect 268402 800 268878 856
rect 269046 800 269614 856
rect 269782 800 270258 856
rect 270426 800 270994 856
rect 271162 800 271638 856
rect 271806 800 272374 856
rect 272542 800 273018 856
rect 273186 800 273754 856
rect 273922 800 274398 856
rect 274566 800 275134 856
rect 275302 800 275778 856
rect 275946 800 276514 856
rect 276682 800 277158 856
rect 277326 800 277894 856
rect 278062 800 278630 856
rect 278798 800 279274 856
rect 279442 800 280010 856
rect 280178 800 280654 856
rect 280822 800 281390 856
rect 281558 800 282034 856
rect 282202 800 282770 856
rect 282938 800 283414 856
rect 283582 800 284150 856
rect 284318 800 284794 856
rect 284962 800 285530 856
rect 285698 800 286174 856
rect 286342 800 286910 856
rect 287078 800 287554 856
rect 287722 800 288290 856
rect 288458 800 288934 856
rect 289102 800 289670 856
rect 289838 800 290406 856
rect 290574 800 291050 856
rect 291218 800 291786 856
rect 291954 800 292430 856
rect 292598 800 293166 856
rect 293334 800 293810 856
rect 293978 800 294546 856
rect 294714 800 295190 856
rect 295358 800 295926 856
rect 296094 800 296570 856
rect 296738 800 297306 856
rect 297474 800 297950 856
rect 298118 800 298686 856
rect 298854 800 299330 856
rect 299498 800 300066 856
rect 300234 800 300710 856
rect 300878 800 301446 856
rect 301614 800 302090 856
rect 302258 800 302826 856
rect 302994 800 303562 856
rect 303730 800 304206 856
rect 304374 800 304942 856
rect 305110 800 305586 856
rect 305754 800 306322 856
rect 306490 800 306966 856
rect 307134 800 307702 856
rect 307870 800 308346 856
rect 308514 800 309082 856
rect 309250 800 309726 856
rect 309894 800 310462 856
rect 310630 800 311106 856
rect 311274 800 311842 856
rect 312010 800 312486 856
rect 312654 800 313222 856
rect 313390 800 313866 856
rect 314034 800 314602 856
rect 314770 800 315338 856
rect 315506 800 315982 856
rect 316150 800 316718 856
rect 316886 800 317362 856
rect 317530 800 318098 856
rect 318266 800 318742 856
rect 318910 800 319478 856
rect 319646 800 320122 856
rect 320290 800 320858 856
rect 321026 800 321502 856
rect 321670 800 322238 856
rect 322406 800 322882 856
rect 323050 800 323618 856
rect 323786 800 324262 856
rect 324430 800 324998 856
rect 325166 800 325642 856
rect 325810 800 326378 856
rect 326546 800 327022 856
rect 327190 800 327758 856
rect 327926 800 328494 856
rect 328662 800 329138 856
rect 329306 800 329874 856
rect 330042 800 330518 856
rect 330686 800 331254 856
rect 331422 800 331898 856
rect 332066 800 332634 856
rect 332802 800 333278 856
rect 333446 800 334014 856
rect 334182 800 334658 856
rect 334826 800 335394 856
rect 335562 800 336038 856
rect 336206 800 336774 856
rect 336942 800 337418 856
rect 337586 800 338154 856
rect 338322 800 338798 856
rect 338966 800 339534 856
<< metal3 >>
rect 339200 170008 340000 170128
<< obsm3 >>
rect 13 170208 339200 337857
rect 13 169928 339120 170208
rect 13 2143 339200 169928
<< metal4 >>
rect 4208 2128 4528 337872
rect 4868 2176 5188 337824
rect 5528 2176 5848 337824
rect 6188 2176 6508 337824
rect 19568 2128 19888 337872
rect 20228 2176 20548 337824
rect 20888 2176 21208 337824
rect 21548 2176 21868 337824
rect 34928 2128 35248 337872
rect 35588 2176 35908 337824
rect 36248 2176 36568 337824
rect 36908 2176 37228 337824
rect 50288 2128 50608 337872
rect 50948 2176 51268 337824
rect 51608 2176 51928 337824
rect 52268 2176 52588 337824
rect 65648 2128 65968 337872
rect 66308 2176 66628 337824
rect 66968 2176 67288 337824
rect 67628 2176 67948 337824
rect 81008 2128 81328 337872
rect 81668 2176 81988 337824
rect 82328 2176 82648 337824
rect 82988 2176 83308 337824
rect 96368 2128 96688 337872
rect 97028 2176 97348 337824
rect 97688 2176 98008 337824
rect 98348 2176 98668 337824
rect 111728 2128 112048 337872
rect 112388 2176 112708 337824
rect 113048 2176 113368 337824
rect 113708 2176 114028 337824
rect 127088 2128 127408 337872
rect 127748 2176 128068 337824
rect 128408 2176 128728 337824
rect 129068 2176 129388 337824
rect 142448 2128 142768 337872
rect 143108 2176 143428 337824
rect 143768 2176 144088 337824
rect 144428 2176 144748 337824
rect 157808 2128 158128 337872
rect 158468 2176 158788 337824
rect 159128 2176 159448 337824
rect 159788 2176 160108 337824
rect 173168 2128 173488 337872
rect 173828 2176 174148 337824
rect 174488 2176 174808 337824
rect 175148 2176 175468 337824
rect 188528 2128 188848 337872
rect 189188 2176 189508 337824
rect 189848 2176 190168 337824
rect 190508 2176 190828 337824
rect 203888 2128 204208 337872
rect 204548 2176 204868 337824
rect 205208 2176 205528 337824
rect 205868 2176 206188 337824
rect 219248 2128 219568 337872
rect 219908 2176 220228 337824
rect 220568 2176 220888 337824
rect 221228 2176 221548 337824
rect 234608 2128 234928 337872
rect 235268 2176 235588 337824
rect 235928 2176 236248 337824
rect 236588 2176 236908 337824
rect 249968 2128 250288 337872
rect 250628 2176 250948 337824
rect 251288 2176 251608 337824
rect 251948 2176 252268 337824
rect 265328 2128 265648 337872
rect 265988 2176 266308 337824
rect 266648 2176 266968 337824
rect 267308 2176 267628 337824
rect 280688 2128 281008 337872
rect 281348 2176 281668 337824
rect 282008 2176 282328 337824
rect 282668 2176 282988 337824
rect 296048 2128 296368 337872
rect 296708 2176 297028 337824
rect 297368 2176 297688 337824
rect 298028 2176 298348 337824
rect 311408 2128 311728 337872
rect 312068 2176 312388 337824
rect 312728 2176 313048 337824
rect 313388 2176 313708 337824
rect 326768 2128 327088 337872
rect 327428 2176 327748 337824
rect 328088 2176 328408 337824
rect 328748 2176 329068 337824
<< labels >>
rlabel metal2 s 1490 339200 1546 340000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 90178 339200 90234 340000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 99010 339200 99066 340000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 107934 339200 107990 340000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 116766 339200 116822 340000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 125598 339200 125654 340000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 134522 339200 134578 340000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 143354 339200 143410 340000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 152278 339200 152334 340000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 161110 339200 161166 340000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 169942 339200 169998 340000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 10322 339200 10378 340000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 178866 339200 178922 340000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 187698 339200 187754 340000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 196622 339200 196678 340000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 205454 339200 205510 340000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 214378 339200 214434 340000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 223210 339200 223266 340000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 232042 339200 232098 340000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 240966 339200 241022 340000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 249798 339200 249854 340000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 258722 339200 258778 340000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 19154 339200 19210 340000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 267554 339200 267610 340000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 276386 339200 276442 340000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 285310 339200 285366 340000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 294142 339200 294198 340000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 303066 339200 303122 340000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 311898 339200 311954 340000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 320822 339200 320878 340000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 329654 339200 329710 340000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 28078 339200 28134 340000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 36910 339200 36966 340000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 45834 339200 45890 340000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 54666 339200 54722 340000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 63498 339200 63554 340000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 72422 339200 72478 340000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 81254 339200 81310 340000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4434 339200 4490 340000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 93122 339200 93178 340000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 101954 339200 102010 340000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 110878 339200 110934 340000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 119710 339200 119766 340000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 128542 339200 128598 340000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 137466 339200 137522 340000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 146298 339200 146354 340000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 155222 339200 155278 340000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 164054 339200 164110 340000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 172978 339200 173034 340000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 13266 339200 13322 340000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 181810 339200 181866 340000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 190642 339200 190698 340000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 199566 339200 199622 340000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 208398 339200 208454 340000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 217322 339200 217378 340000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 226154 339200 226210 340000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 234986 339200 235042 340000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 243910 339200 243966 340000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 252742 339200 252798 340000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 261666 339200 261722 340000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 22098 339200 22154 340000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 270498 339200 270554 340000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 279422 339200 279478 340000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 288254 339200 288310 340000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 297086 339200 297142 340000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 306010 339200 306066 340000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 314842 339200 314898 340000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 323766 339200 323822 340000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 332598 339200 332654 340000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 31022 339200 31078 340000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 39854 339200 39910 340000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 48778 339200 48834 340000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 57610 339200 57666 340000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 66534 339200 66590 340000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 75366 339200 75422 340000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 84198 339200 84254 340000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 7378 339200 7434 340000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 96066 339200 96122 340000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 104898 339200 104954 340000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 113822 339200 113878 340000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 122654 339200 122710 340000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 131578 339200 131634 340000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 140410 339200 140466 340000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 149242 339200 149298 340000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 158166 339200 158222 340000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 166998 339200 167054 340000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 175922 339200 175978 340000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 16210 339200 16266 340000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 184754 339200 184810 340000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 193678 339200 193734 340000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 202510 339200 202566 340000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 211342 339200 211398 340000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 220266 339200 220322 340000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 229098 339200 229154 340000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 238022 339200 238078 340000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 246854 339200 246910 340000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 255686 339200 255742 340000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 264610 339200 264666 340000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 25134 339200 25190 340000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 273442 339200 273498 340000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 282366 339200 282422 340000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 291198 339200 291254 340000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 300122 339200 300178 340000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 308954 339200 309010 340000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 317786 339200 317842 340000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 326710 339200 326766 340000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 335542 339200 335598 340000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 33966 339200 34022 340000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 42798 339200 42854 340000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 51722 339200 51778 340000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 60554 339200 60610 340000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 69478 339200 69534 340000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 78310 339200 78366 340000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 87234 339200 87290 340000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 339200 170008 340000 170128 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 339590 0 339646 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 338486 339200 338542 340000 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 281446 0 281502 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 283470 0 283526 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 285586 0 285642 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 287610 0 287666 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 289726 0 289782 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 291842 0 291898 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 293866 0 293922 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 295982 0 296038 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 298006 0 298062 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 300122 0 300178 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 302146 0 302202 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 304262 0 304318 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 306378 0 306434 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 308402 0 308458 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 310518 0 310574 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 312542 0 312598 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 314658 0 314714 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 316774 0 316830 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 318798 0 318854 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 320914 0 320970 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 322938 0 322994 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 325054 0 325110 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 327078 0 327134 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 329194 0 329250 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 331310 0 331366 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 333334 0 333390 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 335450 0 335506 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 337474 0 337530 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 187882 0 187938 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 189998 0 190054 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 192114 0 192170 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 196254 0 196310 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 198278 0 198334 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 200394 0 200450 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 202510 0 202566 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 204534 0 204590 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 206650 0 206706 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 212814 0 212870 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 214930 0 214986 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 219070 0 219126 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 225326 0 225382 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 229466 0 229522 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 233606 0 233662 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 237746 0 237802 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 239862 0 239918 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 248142 0 248198 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 250258 0 250314 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 252374 0 252430 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 256514 0 256570 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 258538 0 258594 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 260654 0 260710 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 262678 0 262734 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 264794 0 264850 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 266910 0 266966 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 268934 0 268990 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 271050 0 271106 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 273074 0 273130 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 275190 0 275246 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 277214 0 277270 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 279330 0 279386 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 282090 0 282146 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 284206 0 284262 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 286230 0 286286 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 288346 0 288402 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 290462 0 290518 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 292486 0 292542 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 294602 0 294658 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 296626 0 296682 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 298742 0 298798 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 300766 0 300822 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 302882 0 302938 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 304998 0 305054 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 307022 0 307078 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 309138 0 309194 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 311162 0 311218 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 313278 0 313334 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 315394 0 315450 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 317418 0 317474 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 319534 0 319590 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 321558 0 321614 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 323674 0 323730 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 325698 0 325754 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 327814 0 327870 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 329930 0 329986 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 331954 0 332010 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 334070 0 334126 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 336094 0 336150 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 338210 0 338266 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 145010 0 145066 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 153290 0 153346 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 163686 0 163742 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 167826 0 167882 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 171966 0 172022 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 178222 0 178278 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 180338 0 180394 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 182362 0 182418 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 184478 0 184534 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 186502 0 186558 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 188618 0 188674 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 190734 0 190790 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 192758 0 192814 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 196898 0 196954 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 199014 0 199070 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 203154 0 203210 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 205270 0 205326 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 207294 0 207350 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 211434 0 211490 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 213550 0 213606 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 215666 0 215722 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 219806 0 219862 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 221830 0 221886 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 223946 0 224002 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 225970 0 226026 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 228086 0 228142 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 230202 0 230258 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 232226 0 232282 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 234342 0 234398 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 236366 0 236422 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 238482 0 238538 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 240598 0 240654 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 242622 0 242678 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 244738 0 244794 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 246762 0 246818 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 250902 0 250958 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 253018 0 253074 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 255134 0 255190 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 257158 0 257214 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 259274 0 259330 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 261298 0 261354 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 263414 0 263470 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 265530 0 265586 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 267554 0 267610 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 269670 0 269726 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 271694 0 271750 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 273810 0 273866 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 275834 0 275890 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 277950 0 278006 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 280066 0 280122 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 284850 0 284906 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 286966 0 287022 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 288990 0 289046 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 291106 0 291162 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 293222 0 293278 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 295246 0 295302 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 297362 0 297418 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 299386 0 299442 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 301502 0 301558 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 303618 0 303674 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 305642 0 305698 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 307758 0 307814 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 309782 0 309838 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 311898 0 311954 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 313922 0 313978 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 316038 0 316094 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 318154 0 318210 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 320178 0 320234 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 322294 0 322350 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 324318 0 324374 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 326434 0 326490 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 328550 0 328606 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 330574 0 330630 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 332690 0 332746 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 334714 0 334770 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 336830 0 336886 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 338854 0 338910 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 172702 0 172758 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 185122 0 185178 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 201774 0 201830 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 203890 0 203946 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 205914 0 205970 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 210054 0 210110 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 212170 0 212226 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 214194 0 214250 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 216310 0 216366 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 218426 0 218482 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 222566 0 222622 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 224590 0 224646 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 230846 0 230902 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 232962 0 233018 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 234986 0 235042 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 237102 0 237158 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 239126 0 239182 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 247498 0 247554 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 249522 0 249578 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 251638 0 251694 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 253754 0 253810 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 255778 0 255834 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 257894 0 257950 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 259918 0 259974 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 262034 0 262090 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 264058 0 264114 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 266174 0 266230 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 268290 0 268346 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 270314 0 270370 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 272430 0 272486 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 274454 0 274510 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 276570 0 276626 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 278686 0 278742 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 280710 0 280766 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 311408 2128 311728 337872 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 337872 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 337872 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 337872 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 337872 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 337872 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 337872 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 337872 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 337872 6 vccd1
port 616 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 337872 6 vccd1
port 617 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 337872 6 vccd1
port 618 nsew power bidirectional
rlabel metal4 s 326768 2128 327088 337872 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 337872 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 337872 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 337872 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 337872 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 337872 6 vssd1
port 624 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 337872 6 vssd1
port 625 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 337872 6 vssd1
port 626 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 337872 6 vssd1
port 627 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 337872 6 vssd1
port 628 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 337872 6 vssd1
port 629 nsew ground bidirectional
rlabel metal4 s 312068 2176 312388 337824 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 281348 2176 281668 337824 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 250628 2176 250948 337824 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 219908 2176 220228 337824 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 337824 6 vccd2
port 634 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 337824 6 vccd2
port 635 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 337824 6 vccd2
port 636 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 337824 6 vccd2
port 637 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 337824 6 vccd2
port 638 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 337824 6 vccd2
port 639 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 337824 6 vccd2
port 640 nsew power bidirectional
rlabel metal4 s 327428 2176 327748 337824 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 296708 2176 297028 337824 6 vssd2
port 642 nsew ground bidirectional
rlabel metal4 s 265988 2176 266308 337824 6 vssd2
port 643 nsew ground bidirectional
rlabel metal4 s 235268 2176 235588 337824 6 vssd2
port 644 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 337824 6 vssd2
port 645 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 337824 6 vssd2
port 646 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 337824 6 vssd2
port 647 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 337824 6 vssd2
port 648 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 337824 6 vssd2
port 649 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 337824 6 vssd2
port 650 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 337824 6 vssd2
port 651 nsew ground bidirectional
rlabel metal4 s 312728 2176 313048 337824 6 vdda1
port 652 nsew power bidirectional
rlabel metal4 s 282008 2176 282328 337824 6 vdda1
port 653 nsew power bidirectional
rlabel metal4 s 251288 2176 251608 337824 6 vdda1
port 654 nsew power bidirectional
rlabel metal4 s 220568 2176 220888 337824 6 vdda1
port 655 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 337824 6 vdda1
port 656 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 337824 6 vdda1
port 657 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 337824 6 vdda1
port 658 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 337824 6 vdda1
port 659 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 337824 6 vdda1
port 660 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 337824 6 vdda1
port 661 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 337824 6 vdda1
port 662 nsew power bidirectional
rlabel metal4 s 328088 2176 328408 337824 6 vssa1
port 663 nsew ground bidirectional
rlabel metal4 s 297368 2176 297688 337824 6 vssa1
port 664 nsew ground bidirectional
rlabel metal4 s 266648 2176 266968 337824 6 vssa1
port 665 nsew ground bidirectional
rlabel metal4 s 235928 2176 236248 337824 6 vssa1
port 666 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 337824 6 vssa1
port 667 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 337824 6 vssa1
port 668 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 337824 6 vssa1
port 669 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 337824 6 vssa1
port 670 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 337824 6 vssa1
port 671 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 337824 6 vssa1
port 672 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 337824 6 vssa1
port 673 nsew ground bidirectional
rlabel metal4 s 313388 2176 313708 337824 6 vdda2
port 674 nsew power bidirectional
rlabel metal4 s 282668 2176 282988 337824 6 vdda2
port 675 nsew power bidirectional
rlabel metal4 s 251948 2176 252268 337824 6 vdda2
port 676 nsew power bidirectional
rlabel metal4 s 221228 2176 221548 337824 6 vdda2
port 677 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 337824 6 vdda2
port 678 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 337824 6 vdda2
port 679 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 337824 6 vdda2
port 680 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 337824 6 vdda2
port 681 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 337824 6 vdda2
port 682 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 337824 6 vdda2
port 683 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 337824 6 vdda2
port 684 nsew power bidirectional
rlabel metal4 s 328748 2176 329068 337824 6 vssa2
port 685 nsew ground bidirectional
rlabel metal4 s 298028 2176 298348 337824 6 vssa2
port 686 nsew ground bidirectional
rlabel metal4 s 267308 2176 267628 337824 6 vssa2
port 687 nsew ground bidirectional
rlabel metal4 s 236588 2176 236908 337824 6 vssa2
port 688 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 337824 6 vssa2
port 689 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 337824 6 vssa2
port 690 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 337824 6 vssa2
port 691 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 337824 6 vssa2
port 692 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 337824 6 vssa2
port 693 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 337824 6 vssa2
port 694 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 337824 6 vssa2
port 695 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 340000 340000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 129557362
string GDS_START 1235384
<< end >>

